//----------------------------------------------------------------------------------------------------
// This is the top file of the example test for Avalon Streaming BFM user guide
// The Qsys test bench system and the test program are instantiated.
//----------------------------------------------------------------------------------------------------

module top ();
	sonic_application_top_testbench_tb tb();
	test_program pgm();
endmodule
