// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OIrEQNtKhBizaGm0/Sb/8+T0m6tEx3TAuXcVe2H9Q5SrqqCPXVw/N0cwJY+P4war
XD25vasw8BMAG5BhW4qYyVmPp+A5pVffdrpb5XXx03jt/MrHWqgNCMTn7HRipoy8
H3vcWgOLLdBmhIC+JLzRNrq3QRH4sITmcrxV2YpSqOM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16240)
eaMIGo5CYXtus6wxE+3ZtIsNKOFmOViUp6bpLYKJPfwWvJGweSi+vZ9sW8BSayQY
p8c43M/++dnK3C9IlhMDBlfLGisOllde5cf2Do+OHsO2w/bkkVLqRmabkXWyFmlo
vO0mEFSQXX7vXy7Ir90TyBuj1FRH9X+fJ3WjeVSlIotpPQjmsCUCy7IQnPbvRIKy
JM2wz1Xm7/KlNZY+Q/zlV0L9U0otdbgx87Su0PwXKeOcIEP752SxzUQzHETrNtpo
Bkd1wpoz7Rj2nqOiVGyZsVKhqx/fIkSfxcBCJenYK5Bk2ZuQCT/icIUJ/14dEHZS
us1IvjUBh8ahC2ln/6aNmkdiGTpsSQPY2r+h0h2gbVyzqf0EJ7TSBh6JJcLu+sXD
2D9EK+RZskhMXTAbh9DUSM97YwlFqObYpdYYkJ78D9sNV2UtruaVldzG/Ez5YWwe
Z329N5YDJ89/h4s15UJS7amcQ+xw1Wkd+CufY9bc2OVWRWD7/GidEO/zvHnfRkCX
lzxC+ifFTXQjudUU3TueZFKbM+J1dwWtbScfVy6ntjbvRHQYS3DZDeVjZqrAsARc
61IBg5EveUsR3yxjp1JvS7YsfwRNrojF58FutkaQ7H7DXNhMH0QC3/avXwO4eJAS
oH9JsoxiLXxt1I5jTakPGXixbwIoVnokWIsB5CcOuxSYlVwhmqnPV3IXyLCzThDi
iec/0CvD/sn7ePRdLbFZzCotX66nMHupR+2hDot6GZTFZcqKXTudI28PeRCQU1ZM
Vaswl805kK4Y1Q544MLwGPmM+C00/ZM4NGizaWKbZm38mlsQviNSG82MQk5W37G4
KItfLNm0vATCd1N/TuODYhfMs7d30WfP8GPn7DX9bFhE9UC2N3KILnVHJjEo3ooW
wFX6o6xTCrU8bAU9AHAr+kjAfnNAEPnlI298v07UTVKYToX4Rkk1OEBb8OHFkcXZ
fYTi0vl4jdFIwnSlMhsKLxJbbd3X4XKw/rmEXfPyD3nJqn2M079Ipv7fCakoUbj9
K6RYarGeclAJXY9zv8a0eSy4/aRt5cIwxvwb3U4M3vGH7Zxf26POyOWpx64qJPBq
1o4sELSNzDo1iMIl3iUKRo0CJs0eRwTUVoYvhOibaCJb7R5abe4qpM4JbU897d3g
yK7l+Mw1A7t5Y00VmnP1LFwnAG4juz/BNFYceLSLlXd4ZgWKlvzuBOHVcxkwFIaz
QVeFKBUNefgLWXRGE3oyGCdFN5vdJ6Q4nIBBcg/9QFqR3jqNWoinAzrEKLm/jp+H
MrwV8dJ0/60MdrLedGPioNF11/M+SHJCtR8bFu44B2iwI7A2qJrF+MbL1oEWDyoT
gdWlStAUfDru7s+6yJ/NqM51b+vWeBN7/29q2G3gCqGH52QBn66WuOWX3zt3mKDx
m8aJugzvU7ugCJ7xLiIbT8sHtoVLIuCuoyhWYdGyR9IymJswhcyX0KLSifjvWqAS
NwINJV7Y/6Mc8FRRDv0HWHcp+KxB6ehhfaLil+lD6rqCVDcB7DRTg7r/cXZKhVZi
e2rXtAr+LUIdseEE/bAL6kpWd/GVtUyOxvdRV0+0HB/p9g6bILXJYvceevntDu43
30BPTRKg8qj3N2hdEcuw1Sjzxjb62qVhzefRVKZd3Rx7Raxun9m6NJxYpoNwe17y
RvcyOXaKYnuPtnXdP6zJ6DCanBV6utw4PXIipqzXEjX25CpqoTo6IEJHKFwLissz
PaEF/ItanUZR4jO0WPayMeuy8+rqgrYoIt33QtvUVZucEiWLKZpOILuiO+qL34I0
3sdewecyjFK5OasoFqV6t8ds7dlzy6CLw8O4ugp+wfs3xV8QNLJ4XOLSwelLVhRJ
mFW80KlL2IJ9YVqhfPBiLq/b/m5TzkuVq1WyBF/TbPDLk/bNQ/6SgpLkNGsOMdU6
Oe9NVf84/HEni7RXW2WlpeuW0jadSsZPblh7ZbF7ZtLPgfk5/H2oD3ejyMAxlAxf
16naMJ7FYFXGMdGPbXXAeYZmLAzx6EZB4d6tzvP2kPPAQ1tvGg+iI2DOZlWers5M
A4FpVP//lWCFEkWilehv2A7t/DDIIVbs1uDzAIikKfkFJURGP68XYsrL9YlP45DE
KEVYHI69iFBSGHd6HibxAFwY6rCHVK6TxckiI9niFuNapswDC3ppzF7x3nXUtq8Z
rOip3SVGtYcfKr/KWwXT+dDHVc2qC+hJ6oKAbb/7G2RvtjkHAQNp1tGLdxUNwfNK
ZXoV1ktP0PXIpH9Twx3DMsXjJy2XhF3yhJA9F5onYGl8Uco4FEJjZ5L/ghBzrAaQ
cs5sPwgglDKLyq8NPMLTle2OLFbySHsaowY64A+DFnrC8OU89J7Xs2Lk9Z3zA35B
7vljFBQu14FS//4eXWGALhHh0VKk4U5XgdGJislvfRQScOUkrdqzI9pTYHJtg+xo
EYWFdocxCehp+8scXZttWWtb6PcSwpyZqhRAPPW/Sjgv3s5KMfDiI1QPcEgyJ/Lv
qneTRbNvjOG89OrJagvqvCTTpX5VzsEP3ZJchvm2qVHSOsxLWl66DoiBjRfKT6JH
64ARkAUYet7zhDjVYv4XSZhhk9dytexYLE+e60F+2nMYMnWyGNZ/8kxbFvJl9Kf5
NI9OiKArOh+mQaFzKPhaPdL4t9XTYipvUaTGMsfpOASH+1fnJgPmaByOZJQ6KlKy
lY3cdKIjQh6tmMDVp1v7TF5iu9MCc5UcmRSEYpJ2kGsbSxol4kSYl9YcXyql5k3n
/vuaJO1iUsADi/hYhPnwOcDCnQeRgpx6SUNTPLTEVrZ6PimhUQprmFV/wAm7qnBD
sxFakQZrXQA7HBSdMwLA1edbi2O/8cYr8eM1RZrACGScnpfqZHOPrhvH16m9OgCp
2Dg76XnVNtw3awsEwael2n34xgtcoceAG/6XVvgIX8BS5eqOFkPmfkFUjs/enb/F
/TU9l0+ugB/16NvYmw1sf6QIG3ys+564vE+Tw9SQS5nYrQfPJ8M/CHTyx0OtpSRO
tixyL7awnxxiA85GZNA0xAVY7vDFzp97wIFzYIslXNVHERwTXaDDM2pbA/jKD8Ob
cR2pr4jelIQm7ZQHp9PWDuuBRjn0fDUl35fG2Z08Yo8XdbvM0DbGnTIi5bQx8q8J
JGMHARkCP8SYhlMuKqMjAaiNIiWisnIE30FdBzOxaW0Joz4Hvz+78fqX8eA52x6C
VMw5NBDRONnKua9UYdxbfiohhrsHgEhLwR5aLw5CRQ0UbP0lVNjwmRslHzn1lndP
HRNSvy5Hj269sFmpkPszceDH45A2uHlcQxkuTbE5IDjiNDIuKDMc49I+IIMx3lNW
F41XYNx23PQ983Mj5KsuxTpPTDQ+nYDR2zGN+1tTOsTvp1mZ1dYmmd/WxZyjSf6j
KoVyTz+VQG+Qh0+2Yh74r519t5t2wd2IxO/v4qNJYZfxZpp/jKLo2uz2HVF2O9pP
KcRon8VwDprIiyOHDCvxZ2lzEAVTXL3hwpZzoLr0k0NSeQ0yYCoMH/FoiRD8aAVf
Rslb09n0QDqbefxtw1X6hZBWqDaWcPup5WiEmJE1s+LgFYo31A2GOeQRy/41zdxE
vl9z8AQwlAFV9BJeJ3oyld2VemFbXBkDVAlP/BA/Ep3pPZtL8VvSLII1Nt8txlV/
iGkDIZNNlkdyOCPg+pxMCU9u14ioDGJrWGONzrY/R8YOKA+9HM8rBHtAQv241gZW
NO7ugRfv4dNSuwfvTWLpLHIcfm9V4ekPS1jP65fqcRA+5vaQYLC017i4UWTMWzXN
fKDwUFv0xrl/ZrtjfHGaTZYvNO4zGe/82UbXVa9feX4q43dzQC0DATRCEZhV7wQu
bwyYogyrsFwwPrplyrkx7ygDuf/FNss4ObrB2MWtrbgNdD5qL2mjO1HjcM7zuIZC
+SWxKgbc7RhF5ZyeQFQEEN5sympmDGA0VewLXowFwmcZw59BqJ37Np2b7JnLqhKS
JIxaLNJ2zAYZ7TcdjSKhWTsFzG/dmXc7DxVrMNgxNdmlloMS9i/1RBHldVMJbrI4
ZyPBYMFoRE9yfx5PaHqTcloTqMtCo8NKY6uGvNphKK3X0CTFTWJqflqmH1fFoVnj
6U+iyHAXjJMjzBmVIdkuU+WDBflsiZ+NfCK1QxfFiEqAxjGwa2balnlSi8LApevR
ZK6SLhXniYpA/BDmRQYm5lFvBDANHeUe9D8E1b0V7ZjMY9d1uSdsV3HyMYYLD4EG
uh+wQWYrSg7JBAxTI9oQwrGejNcHisQCwDnydVCbVUJjDA9ZBzJhFGMEqv0xz780
y42mg/IkX3z0LZh+y+QLGdP0O0N2C8uoi7WoM24P1w3lZ2iNgUrZbmE1JryZdR0z
3rFwx3bj1ET0wRA0X9hJuQvVPXD8I0uQfxHPVC8pp2jkeyv586d79Qnn0WfSMM0X
VZxIS8FavLlXwpHygtT9BPlW7MuLo9fsgr6ZCMOwf+VuwMksFMY1Q0kEQh4ihOha
Ta20giTbhjgxNJZGy+JvGw1yVv6aCCLLQ8fjiXz97/3jxVsWhkxDExxW7Vr6pSF+
EtqeKCykFBQd9+MG6IvI+wFIw+kRudbk8viqOW7wV/mwKbPmSkJR8b+0P5v0TbJJ
BdoF/dNP7AM0vjxxEJYkV38GkH7ilhj8rtTYR43I8UGjGL0KEkYt6BrtUZIT2D+f
MljP79zXjMA62EtcgIm7F8a7qdS8XJgm3r5k2pS2C6CDuzJa2R36raf3x8WC0JOD
UxI3svyQCQD+PEr38099W7bm/w6Y657JFe3HOvylSKm5IYg3azu8uq6mKIRVeK0R
Qnv59WH56i5N8FyZT+1Gfm12JRtmwyTpKwHpXpb1AP213hMvkYHd1RzG8UraxFZT
rBaXBAtxR/RhN4uLg07fgm81FH4uC1AKWun+0EZ5zPXhpL3Lpk+Ev84g5P/PulEm
pvxVvbKOfdKbQFSNx6pR8T5bu3gcZQqopge9Hw1bZp6cEgRZDQxqkO3dK9GFyvnN
aTjLZNUog4IOGc/MXKP2vHQFMhnptAFJg8MCuuAjQVgavC+4S7G0I7iTiF971OwE
zF6V5boFngtbFfRoiTnu4M0gE1hQMusBBs7wUl35ntlwqm2k6rt0aEbbm8xxMF5n
jOsS7KOsfnU0B/M3wYOA1bIbhO8s1ypV+tWYld8Zsl0HkWi9a9HLq/gI6gTsgOqi
MA3WlmojVBRUZR/OTWTBJcwV9diZexn102owoKb5/c/ma13pPeWhxPeztpFSI313
smhc/Ozen7TpSPVBzNXvFNahv1doDmo/LKjfB6GhNS4nkRxV+bgRu32/cQ0vpcnd
ArDa/Pyov9PcJ9IxhGQUsQsvm6BjYH/4BovC1cC/e2IAM0Vs/fh6/h2lBbwtjas1
cpvw5ixLvjFg1jtBBN8xUIn0aDcfV5c+M6VbnrnVhYf4sH1OAO5z2JrFEy32wSZC
q9wryQwGAnHPWJhOJHI2o5uT7pLfCmIDdJXAct8ZvLsQYB5yiRJ3ARFRe56MQZ+S
fzu9lgRjtvMLRfpZ5ZZVtxmuOMRZUxUP7U/1aVixoH4YRnD8Nwil9h0bBNj6CgKb
OVvDJaaUjFC6me/ThkaZCwcXOhWSFLLbDE3JfviW1uxXp5Cm5mB40YnNiYZZp9KB
93LA2wUg/9vxPG4HPXuexl3uq4zS1bnYIfADq3NC9XK0h+NR48J1xrOcBYz5DAT4
LV+xJMxtyEvk+cYMh6l+WUWsU7Q2pZ1ULKzb0ienRa8HliSXYQ0eD8E0NH06C2ir
fH5rI5iLvhl4w6umjyEKSkHE3LWsr6T/5R/8mkj7T6AApslMAGgZpun8auqyJf9e
voiKYCEOxfVorRRstjSF20eeG/AgH6foUTW2Lj3WztkHXXswPOW3myZBzBvEK08v
RGtSCfE5roSDPXhZPwn6DTuQQ2ta6ltYMXauKVF35DlOcrDSKYPCPoBvKiAmu1MD
R5BRDe2PfZP2ti+lJdu1zhRzL2fXAlMjMS9uEReeHvTZKyLjoikdmuxrk3kBEU6e
fhgYnHvMutillclrETnR4ENidU+MhKP2X7HfcZ8J99acdG0IZk0bk3T9y0Z0Ft2T
Y+uePQ5KWckMJ/DEBVrqPN9DAr2pkxO2mk7fULCtQfVKoYnA9NpryqKVoach4yJi
Mec27JLtc77lO3ptEMxC4wxquKAHmXOOlFbmyd4lryy1w89Z+i1PahAV2jBABK8O
2dRCTiEfpJvkscpgQ332Nkx3Nuu8EMCpCflNOaPLh1s9Zs/X6BOjy8YbVi5KdHNY
f8NzCbD98Fu1q1eBqxqd5uBcHmPjEK4fIAhy5GMhM6ADr6k/QY9aCIrAA7LHWNv2
rzptiyqcx1XFaxgzXy5iwb6+Zjgt9bwV02GQQ25rnOPi3LDR3p7SvWy1jezzkfVS
4vouLoMQKg7paCnZg4aqjryFXmJZPRpuY8nKv1ndAKnLj0SyrJ5vN+6glCPEyHZI
/OjW/H48rOgGmKEiRLkCHDRs8BPDhExsiRM1/gsgFsF83GH/B/tgXGkhA8Fi3G69
y4ZA/Tt5Tk44mMgCNvU3ub9oRMeYFnoz0hblS6kZBExdBJNc/3UOMPwCBCEvamdP
wNHUL7FHic/cG/AzIu89hdeX/LZH9BJLy1+dM0yiPU+WqBm4A9qhB3T1h7Z2tveA
l8wUaNDIZgogvnfHYd5nw9xEIL6b/C+TlSLs2JOGLXuEjZYSviLWIrRNzzpVdzxt
fi9sxzclEMZ+Wk8RruFEHQaKFNagk8zAGAY51+erpbFAHJqABj5WJgVJGNJyq7xm
pjKJOTV94x4GaaeNnvIoZChFQxLBWPm+rw9RLXuiBXouTYNJgmUmEojS+93Zv5pr
MtplfUfH3kCrx/OzPYsLSd76cKQwgR3iTEMZoau+JMPI/md2A3OEIpyUySi9fypv
6LlQViMMk9awm/1ZkrNXfIHC/0LlJnZDF9xqppxAwEyfiT9vzFepRggMzzS2SnUK
2/3y16WUDhlkFFnFilY2LaOLQTZN7qPgNyU//E3s3B5ig00gMojkD3HSNLWaz8Le
q8MSEwR7NYva8vd/pirIVsqL4mA44MoPId8kOLRoZTIgx2FgHzzN4FRXUfCWdvUY
8OqQ6KmBLQjV3AlXqx61q6ffWx4Ua2GVElU3L78WeKqN9mCfRO5JxpUzdcZjybum
PD8TpB9M7cE/o9pNxTN2l8WxuExQqIaTjq3H+6LK5IoPrCFfctc4SwJTbSYTS3FH
JU2qk4pUpJMM/2JxZOFZYYqsClODfigCw6PMo9fomwNFe40TbZWIIRloXRImHBD2
Pc2qskbQWrBGL//dlwFhT0X/I2KNVeMJWlcKtbW9tdi2tLMpmh4jJY8/Z1G94f9u
+11bl4tPD7iTezL3i1JabA2iC2TE69h1Gu4V1SC7iREvvM2EsucOmN0NdZfbKzJe
Sw7FEd4UJ6ew8wtSrtfYYv+6Bmyigb2CpTBOO6rxdqYWV+DxPJ8Df3m1Qu3dCtRc
MrxwSJpP0OoI042tdKOTeBY6NjR2P2VjoIa+3zowhxYjIxI6+n3NNna/0nAMFY3m
fj15U/JsW2sC0tOgq5CmSPGli17F0jjAE2SvYJSVg7+BP1upiMpWdEt8kFX6G9aY
iUKtk7v0L4FBRJDKtBE/j0LlUPm8ZeHNyYSHFzZVVK44agjAMUvmGWnHLtU3FDh0
YUnNjHHTGi5hXmW1zt4awQtAMsqbD7VFGdJfWaOVnSR9suOMp/5hdNF2th68cOAd
l8TKpkpoTx/XC6OrAfUT8mPiUY7jQGz2HPr9Hg/+6ApBX4kge/WARVimEqHiN1mn
sWiwl3BdpQ4faWMxwILzK170tVxbzFDyImOos9n8Fg4ZuSaprIngulkfpjRx/tBS
3tjX2ViGBU4BZxxsCWz6DmhOpOjN1Z85NFhd5CQsmNNCRddkTFF/SBaysWbE9jzk
Vn5tVsAgGZx2ORPyq2635JblczknOqjuDoL9zBgv3s5xCN7NuK4XQlGfXg6q71xX
NTpWtPEss292P1VhHSvNW8TGFvEXwVbeAhjxNLG7sPbtgPDWeTwrXs0CH/lOMn8F
QhBov5szx1tQCvaoa7yPJNquYi817Xu0ldgMm+cLXMAekZUASXYtdB94Q8/P91vf
HpAGSuURrBrzcOIHFnbZiZMlT/+s1LoQIA7xRGpOd1kQ6vzXZikMZDI3yVV5O04w
X+4cgepJ1SiZDTLB/MAITMo6rs5IVOalLIaAjQVPKOGHFuWka3Puyjd6n4w3KSXq
RnuDTLmC7QYQJo/VITtQAfM0YxIR9vdUwPS2uwOu4td+qao10uKNZRTbfnNGalYD
inVS8hXbbocTipa0ZimakG0/O58+ZBQc4c8Hdy0OGPpAvV2S+N3qxHuiEIOry9Hz
mB9hNO9n+Xhz6HvBAYafa33r8H0qQK//NFzhoDEYr12fvtjRAgytbqyXnZBYMFDD
wY0Z2nJxINMp7bG3GsJWPww1/JF+uoFpO66qVjYw9mjiICOm2YZj4ZYfrBGIc7a5
swDQNoI2RplZZzlN4y4iio0fSLz9Tsg2O/4wwcNceIr192IagP6qVTtTsCkQ4ROc
4Q/G9bRKQpRJt85JDEf3RcvVbQ1mOdePQZqLKO1HhN5s4F6p6IQXWX+1CZ45LWAa
3WbXD5PHUO/btch5MAuRm81g0kBFpMKRm4SMTtNowkQ3N/t1hsk9gAhPqWjItFME
GVgkgYxcIbviz0jQiMQPDpChW4tl2djlqPjR4LQOpL2EIdQbvw8CAEGp2/orPwDs
mSBNvgXqYAXYQYasxPlikCNRvCYo3q3eWAN+QV4vl18UXnMgD4Ha0OtrSprUtF7T
4rTFCEWNvW/IkWk8NE4UWGaVVFE3m8X6lzgTb4uAA6MK+s9pCXVa4Af3bXjHei3C
8xGO3+rhyhg0SzwYeTk+a7hxP0ZLAfeHlpyFqkvWa+1nn9wdy+1tND2VHqnvkN6t
cwUwDQpHwak3IDcPMkALahmh5pxrzyeRtAEpYQFOc6XJDaqUGapP+tFjaNVpnB6T
TNxEoYDmZxbmT4/uIaajiSvnu2kVUyqGTYTpifT6EgvSDZBNUGqW2R/8+gAekE+I
cxqzhmxfKry5YqVfLT0h65LnWAql+tDbpGZ1f5PAKn10W//Tg2dSQRSlsEh0fQov
JzIxAxh041uzKx0/SSLsflHlnOuxesIxWQJNDSFpIzmOIDOb0N3PzTpsaIGohY71
UbdHQLG/jkqTOttl30860gQgWu5q+YkWQPCNYLp4xse/DTub+Nv/tZRAnuHdVN4p
bm0a7ABRcvqtVs1ttuIOUHzFDEiNk1tDJ4yS8u9YdgkJTgK0MUTZfOcT+sGYQDBk
OKXHXBYsnWr4NmTjRxZyioeLPb6PlCHt8xov4Illv5ZAlcgMpGeOo5aOVMLGORN+
A8Kfiu1L+Ea+jCr5QEbCVRpVWCzYoqhjm11WJXQigXPXJsTX03dVji2UQZFKT47d
f9/ilDCbrkGUBwP/8iCdQhNKdNvHUziOng2HEFiMirGR6QvOLUgheEkGPhlcF8Y8
iIHiHTj7kvqghl1TT27CqA85VUwZsU9lK9JgeTiYIAGP61Vitk2Ir9uH4xGhfzN8
envVmoYrYQn2mxawt79YoQhH86YOQ0nDzXGWowHZNfqQ3HM/Jx0T1j6Iv3IHpwPH
FZHL6jMJWju3JfzUuTPquzSD9JJZeGEayyZeACjBS6o/u71Ukmj/dEWiWjA8LTz6
ZwJRvesa9fvxYcXfNn8/Wx5uarbfl7JpWrJN6EAuP6awmako70+xsT+l9RXN8+g3
+I7/LMoLD6WaAlgxlsWFh17sc7GSaa3Rt/UP24hpWuBF5ot5C9FPf2apEaCafz0q
X1ljvOaUkaWZYnyToIBovKocNravXXzhAults+4c1wm5FqiW05ErMcZi+r4tzA3x
Oj/iQV50/bILmW3ds5WSX0lkNt3i1rVbhnMhj1wVfEHWDpCZ0Tvu9pOiFl3l9qas
v5d1BZu935Cj+YvZQfhcCeA2zsqcmqZ25/Gz5EKds2yJbPJ9GpSz0MU//x2pYfMK
ejbY61rRd40k/cR5YK/j1nxF9hO9UznyYzbsqwhBtX3TG5uAmitDW3Sz3+u0WtGd
BHfZhDn+q+dJcqubaXshAN3L9oFzZmKrGc4nJvj6/7oIP/LETqQ+kFogHFQO5RtJ
M5X9eGYJkKCdgm51ETsLL9uvAxoFPQ9BStepmtttdlSb6r71LOuUqlOC8NPYdck7
3veuBHe1kjZGGnDSKkAGCKp62zUez3C44uYAPlB7765yXQLcv8KruN+npI1WgdGq
ewdXl9XJBw64JbVzIrwS+wvr2X0lXAH3pYhHiXBdQxGtU0sbW6w6e5MYQXjCoJrq
ptVZQFgJN/izLFaXTL0XAhq02xYFKO3K5s3hqwqUhSUYIkak2aXmVlCRMeXRNwa8
BgpuZmYHiXTh7B8ijAKu6WhKJRje1i5qEZCxeiLcoGRKTyYWaOg3kpyhDmwbU/CS
XTisb9I2iU8YJ8Od8oXe7s4z4SxKcb4mWvTughQhmvwXeqQaOT39SURBo0pbzl+F
jMGZrNXkYsjQdjOTV9FeVHKy1RfqPDOBedRQlz59X4Su0lJTiNwQYqTpiq34h4wV
WHAhiA7Si4jphgxSicbkIKyq2ACFs/6W3/HzN4qJQPV2jB/mw6oMfoban+qcXkfS
FwDeqI1uXWqLZhOIA7dr+VJ1TDEC5PQdy9Mp6VIcLpNvpEROMD6Q8Ze/1YtQFlpn
CoE0wxGgltYM177MyuDqKPqU9W4KoipPhKbc0v7PXLTvZHDCHNzkQGUX+51JWiz+
BpD7Xm95xrdrGSWnWD7u/ZPqeXEeT53DgbAe+hr1+fGMYL2BAKHncrNQQiQVnx0g
81i2PAGNXxxfxyGnBDBXC3krHmH8wljU6zgdqG9UTVy+6WGaWEan27FEHyzv8MdB
VQ58KVJW/EwEBut1ImUhegYUINZEfbOu+vW9zidcyrgLgUC00SVFIQMT/9bC4tKa
kDR5/AFL4gka3+YvknvWNBWhBT40yFfdgnP6/7q8MVmuhVhCWgJ7PAYGV+jo7Nlg
sv2x5Ohpdny2F3AbivonNOhYsnKsd9uRui1nqSovcl4xm92QZfbkJq4wKHVs9gkE
qnkHKPOjuZ2e2YwFg6YLJdj+6sMBUUVWvyMepTdGAEeLDAAJ5QC5oqf1aZEhLx55
RR2h9j4gDeM5VgP+3wjVVjvuNjPnkC1OeNac5ZtqDz3Bt+DY/O7lkb5+ryFwrejN
aTxUZ7wdH2s9gjbGFdeHtPKcDu+2G5wmLgi68ai94lzkpC2QrX46Gf/0WrW0LQAO
DvB7N/QmiD7jjCh0AMUw/yfAVwKqvAU2I3nLnURQWva1C8eMT3G8LDJjiNG3FvJ3
gWwxL6VZRUvBMIjPKl9JbUoRtyyagnp4run3QHqY7GvwQgRQhQJsK44spROkikds
QFxTUA9vo8AKSx2QbxD3sFVRuuOVoq9u3EZZmI6vGFAKxMpkpeVI6rp3WIFM2e+f
Qg02OO4cFbOCeGI6Cx+HmrsCrNGECeQYNt1Z2eKtRCW0V7qVmtAk7tVia+PgtU2H
ePPVZEA63P0HcIZqEyAKPmPooApJC03mmK01BlfB73zvdgLSkwkidx1WfYjdjPhf
ogi79MNKQXhKdFDxShB7uH1s2wZnq37DprrQI5bnfq3AIfMl6GnZCL8z3eANbbNU
UsgjEie7sZ7cTsHUGvFgWKW+zv8ec8m+2EZ+JQg9YofcLTqLSBriH0ZRrVDj3M7Q
eXK2/m+93U6fE6EPUG5xvwrQbAzjwf6tleHXIVMIOKm4skV1dXrn8BIopApcBU5d
kBdkqzLbzg3711C5FhaCUfpxJXOTjseKrEjfpx8655O0sC3BIfIWhQo8BiOk90Ps
Mo/td9jlksebYe8jPXzAZSFno3+pOEyNzhYIhxmsCEH9q39rgL9FrjuxAvr6L5BF
PpyrI7n1NY9FcR7lvzzV6HHtBvFDjc9uhADpPZFCZO0+GfV3PCAcmhEjosGNvwxS
ZhmJeSNOaW1AdoNQ8ReGOiqu0BnLrZEUDaOhReahJTNAs0cCZkCfPMM+UsXNHPnj
ccGpqKddMXPxSgiBPbPzC1+9NZIIJ/abyGmSVxBnvCaMK1ld/eNRJ1y+7Zm0qec1
1WJYe3ASW4tGS7CcZ8xH6BtdFa3UrEpIJaJQu6iWazBzuCJR68nahX3gt1rBcKNE
9IH13LkOqNETZCAzUBlrPvlPq+dRKSdVokhD/LsxiUR2Ul2xNL5y/v0Zez1XF7Xb
VOYCE5IowWHmwoJywMp6GKaFypO1IUArDgTdFgjc3Yobwjto4tnKeU+JJ5kT2q47
Zc9m+yxTSTusshgMGk5TgKj3eEA5GpOXprHNd9aNEaBRlCNQIasUULKpJsuLvfaf
O4VFlPv+P7sAKY2vaHqXxznvWuY4qVZ2neGHrNfeVaAJM63WFZOzAbiqmSCrGThz
FT7IejJ7eIaUQ8Aj3QTv8IBeneSROBxMq1HvLicyrGxjr/4mlLtWey/MKpXbts7d
7OPZxZ0IMcrbrTd6GswwGjy/fUddnL0kzoOl9j4SQ7wolVOY5Fvue0KqCPjBudXg
Dujslc3puVuiBhB3LbnA8jHZGzQnFMSfHRIZLEBRVbxcWagCrQbXZ81/Bf0Dz9XX
LBUFrijWksEEQMWxzmXFKTIJp+A79fZjvgETDTiDCNYOVqUmwA06BLGWwwiDk1xX
vP8fQgeSD7SkGEV3nEZsKYipuHc0QdtZ5JMhKzPkt6RctCEsYqzI4vQ6tF5N+6In
Luf7EZptrcD8xW9i25fmCStAbGIdrzQWKvGpyTo9YX6Mz64HVxd6a48rnyF7PlPi
2DMouvIuyK5GenApM5v9DHvdtHpw+kwaf9lQx0uZyk6VbV8jIOYzK9fRf4I7Whom
iNe+Mzt3uYQT45zFGkNXDrrkQ9va9A1XVzSoMFFoFx5ekrlkzp+7oxxG4/QBpTb7
0aHkKEfEOJ3ljVlsdPuEqu65D+/F9LMRRcONcdZVq73FZhodvxGBoh75fTLjd+df
eWTFBYAkkauNCySSqG6KoP2azRT8Pwm564yRfQSZ4a8A4SHrJ+8lijh5NzIuhix6
WBJpOVS75dm00t95Q99RM8+clNt6razKKgPfqMRqU6ZBvuWN9/BVbvYI6cfrMMcf
NLX/wVP34Jdq3Y3xSwoyYebNbDyahzo5GFS3I+Ki4KbN0iWPc8YMQnEDpLf6WWJK
Xan4eLaJ3nbcf9n6wJMDrf08SUGpFfy7UT6ruRSPK1JjkWpCbSN+Zrs0U62mzCXU
8rF7snMHysR5XjTowkStCPGBq06L8X0BBc9NJ0OOEdtGY9yq/Qq8M2LjngbrNA6E
SVkp4jzENoXzhoEu8lBwQeSaZ4ufcEoyCFiUMBrSGqotnGK6ouUbKxjZ7+xPvDRB
3pFqX4XJ6nlqU0OUQKl3ahIebzUuyvjJ/+NH3td6FCDyLDeAkus/xeRfukVBZ8HE
wnU90GkGTN6OBZzNeFeDfz+4brk5ysBDLvOHyeTiiLgkTNhQ62JE498hv9nAXUD5
D4y6JeYlSU7YC54PFpZV7fiApBex+YpYYcY8wdk9UM8397vJdAz2ng90moGFr3yN
CdrBIjEQ1LlFuGFsfBg8RDLInWJbdXWpf8SYA1dlyzSf5QweEZuUyl8T9QtEP/6K
Dz0gp+75qDHW3WbeKMggcer7iLaun4tZ+qSkGk3F3katXeMzi6wGR65Nwfn0bj4u
lun04hdYZdDAEeeTuv0I07p+sBP+ASeoePKRbgFt18uHH5V972cAFvjbfg7pHGqy
VKccIhVZawaVygeYfc8atzwjFBCZUZzwwkboWLt+g4uN3QTYFwjV9Co1eWqLpyR7
FX2hyChzSeNQRQXhRjlsfFQXyLjNuNP/f0PUTTBvLwc8C9FxlbQkUeVsNF1cI7Fi
7P0amv6MCCGj2Q25squ8IBgxjZ/z6BrM4SPvWMG0VSzk5aF46kHud6L9g5skhUdl
oFOomKo/akLlQq8lb8+HXe8U5n0LxTyjqCjZx+MRj/s2j6T4SwtygsegnP9AXGSK
AxTsurkbHhJuHhTiXjZ4Ne2lV7Dds5EMiq6HfkafhIIJiZyADNzWbtJHHEnVoICN
/BJWBxi6HFbUt7QfhK/4DXskw2GAMSXi82wwcJzqS6b81EOyo7BrKvlt3LC5+P+u
fMp3NBxrPLh736WgMlS2v3kLEJ2U9opr0R/R1QcssdqMAmn8GFFI24fzcp2eTb3w
PyoBJkne9+yo7h2UwBd1dqO/94RXsg5q89YV6DsX47PiGuJelRV38OcfGuvEwXNF
6NgyekhTWCmSQPb9TbnaOpoiafXK7dHWUUkYN6YShMRYvKwVNaZ481IH4G1VGTjW
wvPJjR8bcai4xLBZTfU6tPJ7pugPiq8lh6LQbHZ13tXd0MrWajBzMG6CsX9CFmjz
soW+Kzt8SZs79R2CX+1C/MwxlSVf2iHv79nJrQYeZX+6UmcqAoAA1gy2WGKAy7Na
ImhGl2Zzh0gG9KVg5yBF4wShWEZANrLC87Pr8M+qWxL0rm8edQmHS1nJGNXU6knE
yTO585DHNd0tQveqaElKoaXGQMOvQAdOANWf6/hoIe2hrfi+xn+6TmbmFA30+RD4
AEfhfzXcYkhflGHVsv4hAfC2vFUSlCgBsBqOJr2YoYHYBW1f/wmaSX0ySQ3YLIEA
4QP+IF+t7OA2uaZUb2nyHYGT7fDiCmT3rOH67Ozje0+eDqCiFPCMGxQzqNp3xvij
YsRo6ZMmmQpKkC7EhmvNdBej30qk6UZjxmLoC1wL+9bRDErNxpBJLCiRkh1ydSAz
dmoZNivOWUfYvkZCiV867Ic/dvaIfojUXYQK5o8K9RYDWwu/CeWCE0q39kgY6hZV
14GOHWSzdSYxOOeWGnrwA9p75iPqhuiQP/LdZUGQpkrmacngQghM+fzYpa23dBRl
wEhNRS+Xw1sONmattu5e6m6xZc+k3oL0GLQLTYFULLLk4Lgn19IGEIXorv7cDhWK
YSf1YDw4ck50AUEfVr6S0YoeG1b15GjLcLNpg2OT8VlixmiIhaxxsIXbg/2LBPME
vGfnbpOQYHe9HWRjLl2UX/uq+IJAe+Bt/ES0/Xoy8+r51L4PyOF67PjIaSHZGPQG
ZhTpzrXGQoBC1F0H0YOs8dLSY7NS30uQkOJqCxGAGZzn5MHPtU3Ach5UkuxRH4Yj
26HRoeZzIlPDiiNih2jjiecwzlIleX/s4NRtY8m/duuzIaiOrXFrhCdO8XwKtQ6D
mfi/L89Y5G1DyfqUVc1giCjLXIGR16DKxbtr8aj3twX7eVfTl4Tq9dHNysZFb20B
Gj/8Y4+1kOIopBobRNQeJjhmZnIZQREW5zhrQdCVoMqx6xXoevrvFL1S+2g9mYWo
k3JUKX7n8TcORZGKVb6oCgos5Z/X8r4cBpAnlOvVfAntT1vn8Q0CvMZqjKsreiep
nMP4lx/ZUkvyzmpOfGHhDw7ziYxVdhdM8IoJ5//+6HCz4GSiKaDGsEj1zAePZl3T
RHL0fjoZS/lVDNk82I+xlZROQW4Xf1uZrnTTYzm/3+v6OB4XcrFarpR2I+JKQT65
qrH/g8wVVbi67gglG7xPqB4uHm2l5odmEHg0edt9aB9zNcjtcTk8vJ7uEfjUgtxp
lQ+vQHGoOIBGCJHhxpZfnebCOMeN910bU9Ubd/200QtQO2B4JJL2j1CFcBatutpH
uUQyZWreIlX4pt/LjTKmH4TTq56Ty6h8CqMYfqnUdE0dvqNubYLkVuBxWzj0rcdX
y7ozt9fYmxWbGy5YVm+jvhlA3nYktQbhXII37JFyGtjtHVxFMIIO20F3L10uItav
eUPATnyG9QhtDvTp00KK6NALYld/Ib4Z9w8LMyCBD5s7qQr1kw+bsr5fn07Wq3a6
5XwjawN9mTJ9OVbG9Ay1kfhAFbk4vqGolcFxzxmYc0jhz5Ghbml3IgdUFFbypi8s
WFNYPHoJkLED+axe0Sm4HoJDxhJVuCSHI+Wyc+ILr8OdinEQD+AKv/iDjYteKVc8
y64m1ItWIN3beUzxouN+3VzOh0qppIlMiG2YnQ/6mrLyrDVDNywqC+ih84s1vR37
ntg9l0f4Hfi589KsRxHLxUpEPfa7i3gkK9l+fP5Gkfr2Y5FeC32LyKbhIsGRI+az
0j5hekceFxPOWMdLq4nLFDfz9eNxvHzqLKBuyV84H/+6a2ujAuZS1kvowp7iyjn4
BSF2qia3hYvB+5Rkn3SBRQ1yyvANbHT5kg1Q4l2OqttnTUj+Zfxertt3s6+UD/IA
KUX9W8ngbX8b0bpQFWvBnPb+38nn4zvgW0zZP7Wkbexd0L8jTILZnLeFFPhQgffb
meONk4JN0TAU0IRm8+TPCwrs31gDNn6fWY00Ur+0VrHhLvakj1/GGznzWQQPloet
+Fc+OZjXRXc3/YceolStfumcf4WhdAT1UYnqGp1PoHoXC8e5qT95JYE925wLGzB8
XxDrRP7MOhOO8X87b9+kRGFDqnqlBryyjg1MeMX0YIaHbsnIe6iUiRJRObikAueu
1h0uqqylPCkfrBXxIxn+SZ53WRI99r2rJftbdzqiY35ct6GcUw820y1eY4w4g1Mf
s7quCqygpq0vDzxSz8bHmzu2oyu2sG5qnkW72XrDdBH/lH21Mlk/LQ2POjY4Y9Y+
n2zJwqWXo8SWzpfrqVAJSqmXrWqKXNMd/sI+jRFuoL55E0rKnB0mg73YGRBF2uae
p7Or3yIq3+HFLDjZ2tEGLauvp4hCoQXjwM1E6JEGROH7Gwl8sWnYkA/cPEpoB13m
/e0rGzZw1mmLpk7N1yDBE175tmoTU8RFeao2gpQjk3jBn1FMiqewifKkCHSIoCWW
7C3QkPMetUplXOnpqW1kaEa6g4Yv9rxforOjJ8JXynqGQfN6XGYVNFNHvd/ifgAz
dhhkKYWY0Vnf+AUgY2Cvj1LSNMCM4ya00W+e5ibdKSL+Xllu++Y2l2zKLFOPMydW
JynqEqL2vSbJddSngq37MERE4nDnMtar5gFuELV078Vdak7VvLOouy07u3cnzVYR
72lgWCt8rf8Thu0sY4T1OseLBlYASiI4uJDj6JA03ewF+uIZxR1TkyeCpaHbIXNk
PuOJEy2tOl4yisDRFZCRtUiIwxqnu5PqbVVZ9pFlfPacziUoDbWUIiP5EQTW/otA
k9gv0PATIF95Tb8EtwNAToyiAB44qt4z2IP4GQc3HfrhcdIsy0l743kD3aaHadeX
fmdBn2dWAVgNuvdwF+4p7BdECMGdykTqYT3diqdViDhW6xANgpluz6z+Hofpr4ZB
Is3SrVPxUvlocvMJwRAeoJoy4QbWBYXjxin8P7AX3YSjLoULX/+M1nn6QT/8Tli/
Ba3nAARngp4lN4YIExBV8rLBGFkh2/u4xUllkMQ9X+WhRfqzUeo1DB56ckUSmP8N
Fir+mNx2epbvmTE1x/n1VEWOyPch4PXBdQ4eAr04dHdfcKImpTAe3YD+lEqws6nS
X30o5/ZEXIcbdZ7uaB75Zg2zzFOTND39NrIxO3les2Gj1tcX64IDSgSapHrZGJEH
IYRnFBmQvLgsIHd0XnBxPM9n1P29M8xZNDxOSYOLnGXDIA9c1aZGuuvzdWmO1Ve0
o/tbKyp+Swvt1V1UzCmcJadQnQ/7HsrUCuGobuRY/9fuZbFCXr0XN+YUQG1ZqoTM
iKMYqAG+kJCKvpUrl2ktUDRKOUr+LiTm/pYa/ZiuDEX45CIvH82neRABLEZVJHFW
vAn/o5vOuRMZZNLXLIaRwniymKTppL2KYmpnIDDlIhzOZA78BS71BrZhoXumBptm
BAjfcQWc/oy804+alUWAv6Lf1OBPAqkNBwc6pnz/9UUxsUkY6hQgmI0bv8rgrifn
98thgjhbSe56z4VVgQVM2nc7QVs+5ZSiDRIL5n/rznuHWo9Rqg7+vyEcEG1H/pUa
T+XRuX08Jq6eXWCvqHTMvaqazNRKOYs4IGrkhNmlGDa8JWWkx2hK9k8I7mTQmvaK
7wnDHIKhUQh/E4RRMrpSNWIa+rrMKkrv4If0Zjf3qMrNjWyFJcFvYHmFAK7WhpbC
QYgi9qhNbflIp4V6eVPpp5j/dd+inbqKLB8yBGXLriaIKYpMDH6guvc+6FMX/hdf
Os8cg7Fj+Xuuo30vAYOweGajSVClU3ZiLSbynN1NQo8pBYCSE3qxkMLv2Vmnd6GL
Zxk4+EycusX3VdX7/TANmvF3AQRrYhdqknie1+MMvPTZ6nXYNXmlUhTF7S/JLIdV
IRYmoYbNFsHO9iMp4s/0NOw1HOgJSJwIwCElU6qtqOn/KAOiW4L2i50DFYD4g3Vg
x4ZLjZoGSlV8Qhq/qUa/HR/FL258ltSBOCPiR9vcRWv5AQAY/tFS8GGhVo8ophXc
DV7cu6NHsxbBHRlT9c8h30VofQ/zFOK/LElzrKpJeUYUtjDULR+MpCgNOL7emnHd
hDYUgwd9NLi3SkcrhNdzcIe3TB1AdZC2iCyCi91nSorPAsE2CyS/LQKcqQ9G0JER
QzUq+4Ye9Rd2f929UPVPAM+H0CLYXcwYxcqjRcvPjNBpOT+CdbzGiAemAFnZ4QIr
WVF1qypzO4MyqGjf2nvzFFnJ+oYErvvfmffCQtm+bwcBt4pUKZ2T4AD2hUd4KPeZ
s8fscTU2RDOkKpVqqdyzLqbdv/KIKGxWvtGeWbv0BpKEomqwwyahrBB7LsPDnhZ3
s977RO1QSan+rdPGQif2BkKNmVJcjGXLjjeuCcNduHT3knQ2MhsjIyDX30bF9UtV
59tNeU76HFPzdM7aKBdptx/s4qDJfAi7Nh7NFAVOdcyEwhRu65r0VJLNHYxTs18c
UmnpjVja3WeldM6miZkHGXhannNHsg9XiR5cFCCs6v1FmyutWfAWlJ/3o/0FcMOo
fP/u8N50KvF6Gum3Ug7HKXK+gdJnPgyQRJHOhS0Ru9mVzdOM9u9t2kqL3OTZ7cKN
DR/NQJKoiBJwmMx+DrsI1NfU+6OaGJhlQQwH8dwFMqerveRXD10vnDbhnWppn/UV
i3shDWTsx+uTA8o6Ic4WJqIccBv7CHSyb7f52Nt/L0+ZBPbqmupN6oLg5MGBmEuC
3/hU70RGuuJLEeZh84Qp1/KfQxVTwEay2+Mc7aJRbZgY2ieaR7SqXLgBtX9Mn5SL
2cedoF5SYjTgp+mfDqO3mxZAZljoF4DHoEAc61NBfh58KOkLE8Y4Fpik3OXKNJ9E
16wqc16vAQ5xNCOxkQN/vsJ8xDqPecAPUk86+7wXE8Dj7mV7QMe7CQ6Js3hxpsXa
EWXyIca9G+MZDc9zi46dPkQ+lo1yWs0G5eRRHHxIiQq1XFAHQT+pS+rQXomMBVs3
7FOti+z09o4k+PfatijtCmmobjdKn3MJvPvZMts1CpkuxW8LBb5gqg0yuMV/tcU+
kCfYWcJ74FcAGLc94iraYT3tA9ll/1G6EMHPOfYyPWVbSQ1/KqpSf+A9ojRIzEtw
sbVqLrCAdpmxlmcheglehQ84tafmf8hqLRw2ZDUCdCy5j/X3ZnAHoCAJhl5AkncF
jadIAYLdpX88w/IocBIgSqbF6qZzq1i+hiCRPQhd+uNZSqnpj+xkbxfOyP7AJVyD
2jgKW2zjJav6vTA+ShSDmMpFbMkrZdhnPLIX+AX4vBA/Hu3XX/MgJpbYNulGaIbJ
qkoTiH1eeIzEi1sY9TGnpNz9no1d625wibTMToz4GqW0+Ex+PMtcCXQ1N2CJKG6O
ALKN7astQjSPbfLLtG1my+I3ZjlBriEi5ly0m84B2SRkW9bzlt1r8z1UmONym5E5
+M++FkzxoLHoZiOYEJ4Oi5ZlIiQOUxSCYrUzzJ1b+H316iOypfeZ1iIk7U3JOUbG
/cs91YRfCp8SGVl4JHFumzrScP0nDD549BLQ5UbU+0GueGNkrmtvqv/LI7xLY9X+
m/dO/KAu1CpQFi0x2NHLPOByyHRRhBI4enPhRyKVIl4MxnZkB3KUXeKwkk1xNiYS
7gepUAuCX+JCmDb9VSLAQrW7fHJwrcEcE3G8GIad+cyAKhd/nqm/1f9DEepehvrz
siwHJ64mYijKOGXGaKIEThreK48PzLXvBoJ77Lt/n4m/p7lJSQJCFC6fmgo0+XEj
hAtRE7EiD8XKJg3SCWdWxKj3heyoNge0GHl+ATmcktgw/Y0Cj9r2IkPgchCTBMB9
JS6YUOMmZ0BUf13Xj+yPrIjETd0URHF6rvCiikDJU14KUaaodH/SoHIumV2NYCXz
QR9pFxgys1JpPc31kSMcxqBYLNISUKC17O6MRUp5hbvKayG/NpS26iOyAGfxa38A
xkLvpP6uzKFxYt9phEmdh1PCQNwyTnYZQqeYVIVXh4oAD1ShtzJmESL4oJk8Qmql
l5GmP139OTOx5Bm3KbLDymMhJKiFfZjjAruMuoCHVZJv2Y/g9RhK8gwN2vcERWna
ldzKnDHfNOuuFPmmU4RnFr20zpXRke0NZ/e+p7IkeZ/AO+KEUdjzHBKQasGUVFDD
orwgYy26CJXJwHX72+rPcpdLhfayGWOnKPzs2siU8NnjPtBJIqqsEmyAIs1LXt60
ZyhryAUjGyc1ye2aVuCJyvYuR+JQjjwhgCHE3gmlu12kj9H3ErgYBv1EL+90btV7
S/e3/OYBWp4iISqeUS/E2H5MYx3T4lDsWk0uqX4N1v4PvfC/VBjr6qzeviAB380S
7+N1mJl/GvKyGOJT2RTjp4nh7J1i3gFmfSZO2ODzIQNrLSthHD6t0JMcoYiy+hrj
XjYYxzH/mmktf+9J3JGXYo8iH6SlnMx1tSeDCVhb5cjgZAVwMSTubGQnOxONLIBY
sTi62eiY4OIWL8Ei/FXG0bRAJCN0HqWVy9uA16dNVN9Nt+PxzaevgoYqrvPS5cUg
6CcGiQNrsxdNORl2RwyiosE37BapourVFwhtPPEQMI1ajAuL14+98SlXucVfbpJD
/K9TP6mnIOEvQ5yOS3xP2kqfN/ThMNw08NrmCYi3eIgp7OceYIw2GbkxkabJfXq/
dAiuYaD2XI5Wp7/C4wexvqsMF2qh0aBGsyGBCC0mNQrGiKJ+T0yFK3tZpvv41a9M
/v0S9N7JYl1qnVl+K2nIREs+J6ror/4DKv8cE6Huvk2vkyOi+Q3S9QJ4zMaIjrsA
OrCQ8F1s/tuP4twJioY8y+fFyOeFguIPZoYzFrRvzWGgBVHZW8qf/zp1x8jEFpzG
z2w9XMq0MwKtF1Q3XEhSJOVT+peA40x/1N9w1qC7hSga/oKyN3dXixk+h9s1YiJj
tx2WMvTtosYkk+pCOHL3Ai/g/gmWbvDy4pP5BDb+lop5T2gCHo6Lvi4Gv9Uv2n/E
NLpF7v5DKXYCMmxUpYdcP0f57oSG2W5Xt6H7TKwWcqD6p1wzAqKle/gzAOGBJzmG
7khGLNbyt/1I2sotwzgo/Uo5DGhRdtZcEx1B31Y/1UJhSUlxrcmSeV7BR5P7tE4+
+CR/+klOUEqYZKyZVR7+j77FO/g1L2kXgcuTRIW44h5/kLrm/gLkXgJm8+kaAr5w
RvrOC1lIpg6prrclgIJzM/pDsOPl1101pWhXkAPI8InfJ7qoD6TGbn0rTPrvV14Q
rPWv+Uib1hMUE5r81Aw7FQ==
`pragma protect end_protected
