// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aWnAfWc72lPTphQdylCTgFMVutmcKXlZmNGIk/S8rnq2RfEOF267hp70EG+oMIQI
ks/7av5V/lj2jDm/23E9Cjo0THH411/lZJlRYXo7i4q3aETTW+IpVmmEKqus1Ax0
ZUvHdZrUqwweN8JJjGID7Q37wdkKeNBizpUwlCvkK/k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6576)
S1cyQ3poYAlFl6JKwy85tluzojTlJKEFW5/agENvCmqSUqQVCIImQu+I0kACTpPh
mnULHCbHXLfnsklWKape6CrxOED3IEjn8sczOoiVLIKHh0MT1iiRBDYGN6Aawe9R
YT23/PC5CsudWJxXLNyFAhlXx3GH9s+sjwWHyzRt4o8MYEO7dw5wPzlb7YfHt5Tj
OppnMY53ZdsKaT2duU+6N8ZM1D3OzY7frYEcPPZMHsxTggis5FZsE8bC5VHULfIF
BzRVnmpdmAJrq0LZXSrTXNVKuD+id7piB86ajTq/4FZxHG1YtUQAXn8hrO+j8edm
EXI55YMy3YVzpl5624mA7gUhIcSa+FTFJJcV/HmhsbpOt8sHhzVUulYf827rp+7r
SEDwuODt7O8tUK06teC6+P5RFd6/UJxHCNsJSYuoepSyGneKtY6bd89G0TuHyI4J
ga/SlQCrpHceL0oRxB8CdBsC3DhI4ZWRfk8r2l+LLohw9vnSZiXN3zg/+OLNyjBG
AhE+xU2V8QLXrTAe9VlujlDMdgfVbqXEvcMGOxOzoSYGwKXcGI16MCSdl8hnOXiU
87yF1TXBYLeTEL/bmZHeSK2h4LsHnoVLCodYUp277CXzp/pFQ0oborzSSPBa0vZ8
9FfVLi+CU76gJJfMldfBwmflwkzejhWvsV71KXO2tMVmwAQyODTHI00v8jCMM5G/
oYD31ulZaCYGBJvlk8DZ96HxSKspKr7FRTP72P/emXcrQRvr97Yz0zM3W+LAR0hu
3try0O0RLzX7Inn9iuQnowpRtuHd8KNTvnYB6VYNcv2aVuaXdq8YE4Nxgqpr4RKg
97eUdkd6e+VlUqFY63ukpmj5Qf9XrhHfQAE6M3DFAIikiSpHCoDe0Zp3IwA+itY1
XdLJs4q0Ui6QS8WjKPAr46xx10mOo13iH114vd/9genHzZRGdzMfx08Ncivawn1P
jB7TW3Nc0oNMDz+V6Ob/5wTynezFcnKTjrFv1unbaxzpSCGO2sDqIpDXJJGuyedS
ozZtQUBQl+I6xPCy2MdDlmpzvuD+6KUnFAUaplbrY2y40bHPY/Vfz2FK8IiCSpJo
NsFcbRV42LjlzXBghwNll3+Ny5ZF94nJ7Z5mJpSjF9IT+mccC5Gbm98DGGdioS9s
Wb9QO3ojUT0qT2k7D2GWbEJCOFV9YEOqivP0C2wuRSDvOeLpCzQrrv8j0CvirXv8
4Zgptip5wXF70CbHFM8kjV+ZH13c/Rj8PLOGx/JqKAsecEkHsKAk8voqZ5dQ9aCd
orYB9+7criyLTSgSQtKXBGmsDoC89Ny3iGi0c8nqU0AlkT0uSMJXL7FtYDNEL+nw
OddeEzN3UC76tp3f/kL9/jW9Vzv1zT8wl6mPykIiDsT547o3KX9OtEdHNYKgY2P5
6oo6XOjCp9vipw3rSArIchgc/wD4CZKBQmApgJikEIus95J41iMKIF2e5+7/gECZ
cNG69I/Shm9AUWx1bj9TRnuFEf5B8vgEX1y5aG+sf8M1Fn2xlDkvW6KnvT1Yg9+i
t6+4/iTsxEjQ5vXHVgp9cCMVaudyoHQ7m3LwaBIQXrL7RktlzLsM4NJDyvedlvTG
WRHQO3gIbmwULtWDLlcGUkXIzp73pWhA1TQmIoe6uvNmS+sXVFb3i4VP2yvqQ7BF
NzSY3sXiEN6l6mt4BzhAVh20dUfggh+TRScJNXVgzqEm0FCfw9jlNJhZATUIQ5GS
FlWy/qIHRBd/jeyx8GALxf+yBBOYd+JAPdwqy0/fMWmgWGevV7IRLzjY5IiVk1dB
UIidNuSKkfz+R7WxicIkTafrsXawuSuTDW3pxVO9lC+5oAc6+tLZeebH72CAq42C
OHQWq6Kxova1E+6BC7qW8hoWHnT+wwpRXpyCoqDNwW6mqYqxyawuRsZPT2Yw79QF
oTmzb1zBkoNNt7UGlEE/YxWLPg8NRKbS3eZSND4aYz+ULp++g+m4fOaXCXgXg0kU
QLX7lOcJMTUU/iraU+eu5cV5KJQ4zTgaOatAq1411XVcbvCN5Uzb9Y+QcaAJTkPS
9UFJSD0kzA3LcFdudl7rFLsf/OqZ+ScUMysUBedPYuJonkH9Om0toS86MMTJkRXr
J81m8deGdagY3YyC4Zl1+pEkXbePRhvBtaUKpcA3IGNVBlheGLwv+5S4xuAIVjTv
kTAWmSv9m7CEXCgRtq8yaQ/OZwBmJNyu67hsrYAo6mpQUrD0Pen4KFFRphgBjNDJ
nhM7+VvrJLt/yz+KM+4sW7ivlfHhlgFIYCk8m2nciPAOqUsU/rJa6H41K6WHHclQ
PuReNcvqvUneTZZRxHc7k/xEQhFsixBra4WZNzPyALHAKo2KnGGWPLaKB78+Ndyt
KlYhQftl8rEZZLjrMOFkp3b/HsJ85AQzQWgZzbQJ2VjA1wkPRRcAG+C35Kb7KctA
fCBYitb9T+YizJ4D7jfoIVrH3yQ1w3ES4GNNWC8OPB8h+/+hVc8RP8TWqKmYVYEG
VTu+r8lOpoxFiI7RPiq1lI315r2oQ/6u8TuEzizNIgjS7fuddXufD6ns1K3M3a8V
3IqANIHcZLn2vuNdXfEoOlrxpIk4G1jkDEw3ElmTfMRahNx3B1RGL7/q4GZJpiXR
sSDJ7sMuya3e/Krc4HRoJ7chE50APDhtGMSC1+Jry9B9KEP8qfe00m3E1Gb9lJ+e
jDOeDYb38OLce20+Y3kHjgyZQVNyAFP7LdKwG5qBi8Vzs4THsbPXUqYMN8WkXO04
BL05Ybgqzo3yeZqD+V4fMAQZ3GBWJu6jijttZBlFaTkR9JvidzKd89dWG3i6TaFl
Ofy0zVLtODrWjoCkyqva9qnsItLXCAa1tLZwBYk8t3I/gqLPolY8lwbs+iHUS0nR
ieEX0Vy++xuAgLcT7D8tGpio888d4MPYzHNbz/cYIatKtmw3EsXtq4MlXave1EIH
0zkZug27mBqGVefgcgCZqTcd7+uQZsm1l0eyMQryeiN0/FjpDteHsGeMWnwTQN33
MBFS12voFQKejZ1g1sWrVH/CO3HKDE2BGMLn9ys3q6BIdPqXeSfSmqhw+THckAij
wP9voPdSk1P0npXoDVqo9btRfV60vXaDlM7N5H19zyk9eKG4Hcow86qhpYdlvmrK
x0TIZirV4UhyRfT/jgPq0gpiON2XOndSvJnLxUxMuAGM56BRhdXefPaNtYDpzolr
nk2dhpZoh5am0tlHIa3twIqentCFNzY42l97oE27urIb73Hyo56AuyG10E1+PplH
S1qAdkluu+XkPLOFLeAwbxLA7BGhwvbesI80jTMGshhIin6PwpNJeyIxyc5f7sYQ
lc+yWZOmR9ZBBgUcJ1o40J9N2l7HDDCqUnA1ibJk9OArbSfNw7ezMWkHtCg7MH0G
uo33jcC/8lBpiQ8Nd1Jn8OH2JwCWUCAQZnQexGF9vwDxr4frIxhVo19yQbuZFAyW
5zn0n85IEpVEwPNeaXpPAVNZTPGnKRkQyzrgrUqlr7G0EL+Rstz7jFvHTWOWFDk2
2cTxQIS1ckm9totvC3K65fVNSHunFJa0hsgYpGQqgHDEVd+HoLC6RlbOA7z1tlOV
HdSB0lf1CHAsm4LX3vbJqtzssDKOuL6kK/mw01Ix7IW1ODW6lNuVnzG0TXkgCdY0
UtQB9zwIj8tctHMplsSSxTdZrFPiAGUxM+kjb4ikds0rLIzEmkMMTJG3tCFku1jy
f9ahdzu8/UuNzwuegXnpemIWX3I9h/hhBHFcJgzzHqD4DWOihQ5YUVjDc2W/IEWk
xDtwX8FxP1cKgUCfpaOdqcXb47cZGBbalp89Rs/VmiKV4m71+vGG0bpqJr3aQ5eL
wbxZFi/uLwvLc0rce+JqOknL2kpzabJOn6MLAW0xx1w9KaO5oMuRdPg8fmoZMVqH
FrvxUmeDlclHdQG/NR0On1cgAy2Q3sj5Yz5TVYI2E5s0mIFfU7soV/Lu+mKU6C5C
0M4LdPEODNznAHB1F6cj+Nqv+5ECvAe5oPyeNNIKeo1fo3zUX6lsdkt0ClDLj8tz
0BMfffE7gqIIWjSrozS4Zwb3n6W5bD0iEERkKt55RbNOVJjOG1wmR+zCgRCNz+ml
Wbj/BXnlLPoADe7G1U49qJNelbbRtSETdFSN4DkfwwWcbuke+8ZUGHJuB6LRe2RB
eABNypGVYnAkbVkYNZppKPgnvuROkzlBhwPBmQKhWPkyxq4vy8H5Y5gOaiUBd6kP
EGZi5P/+jmy85LbBJQNPR5BjhG6xtmwzHJQke6/JLj6Qe39yFJCiVDWnO3BV0rGx
0YZ8wAEC7W/eudJFzISVwtTBIMvptPUBvTnXi2hZvygas0/ErrZhfwQKWx1f2C1G
3FpQ1L0OzpI5jZCqd0j3Urss61m0lbF0cbQ+H8YPyN6C7kiBrTr+rvQCMLEqu/go
stb+m8jNn2hDH/BV+j50K557cTRFz4vDELrK0+qgY4/VpfyR+3X5kvvSGiUQhqZx
Xu6RxdY3y9cAt4OYsX0mWUjFPQnXKjCNVIA0AscjAmPpGsXOONbKvokLEvN5wvlR
sZkY1Ok0nlsA7zlynEUVe2VFEgacXEdp8rVRJGMJ+7EMM+QRrI+LwEVMhiEON0Ji
pkgjF5Pp/cElInKkjUDBXqZvOJo0NiX8tTNDbluBTF+Jsm/t6M6/6JrJogvtHt4p
pkvLO6XRv8Kw7QlqFdvhoXQG7O6tHiadvCWL6kDWSfi6k2XHGh9+lkjSWjB6Jgzq
k/d+Rj7kAsN6HGN5nqCm3cLwh/wn3zE5ijiowT2ikglERONrY27u/Pq/GybFXpl6
oRzSFOpS6Sv3hAwLQhrlkqmc3VySy5o+4g/fNY1imXolnWl3LzUduNW8SUUUpPHP
zc7x0+rC2kfLpd6tOGR3LQfyM7uGWsgtT4n5+z/3cgWVQTaTSnGL+f0Sm+2Oc+q2
BZrAK2V3ejJEl0h/9aRGoZMEk2+rQnIBbwmxqmjXkmIDNlzhmC8Jsu2EN3/iEufr
5YVhBcLA/iRdjVKdSEix8OA5B/DIkNu10Pp0PqpGXMZNCTCqjFyKIsTeES6C0L+h
OsSXVtKifmk8wFmlJ/z5kDkM+PesdvQKJUNyS+u3uJl8F2lV9T1E/mv5KeXpt1tU
KcY5fA+JZbTAZlTpn86w+PjAEOpPYSMGeKBBNRXxocG+Wcf8as+lPOzmTwwMEoUm
i2SMUZckV1Htlbbh3XIDD9bJ/gqM2mCr3dPIcQoBtjrwtZGLwThgdxWxyixNUpaS
5SXOulNnPLU25a20t9fkICa5TrsL/99+BeCe/aichXi3vBWOv3jbP7LUXZk5e+WF
McMzFoFfksK/HijpNSzP40L23pbo7C8b7WvAiLSTdkFtwDVKs2lIu5ASvWJ9I3Ru
7ORt5I0yMeXC1fc/lXsuMSWAXzgAmWdiPpBaSzMGfFj1sFgDKtZ1qUUJY6DVVkWu
/PKm3u/mvDYGUHVXJPl5DoV++W1AxzpZxk6uP+HeoXA1xZYv2tjxOGw39fo/3uzK
dGvUIq1Hm43gkrjnlVwgZcDqYV7qUvJRq9UZbnbfaWBfhrDxL5I75CVAMMVrvYnm
pmzhnxFXejFS/mkqKyiGBImq4UPF+oEHon2EEm9cMIIpco+3Wz6lL3cI5dX7IvdY
nVliOZYQPSIb1N+LBza3BVJ6KpFftna8SqGcMbFSGF3EH07Ym37UrJcxFGXPjnun
OXw+9P74/ZQBM4jrmN6L5XAKDoFjIhk/aUNBwszzuoWLFUjlarjmAtH1AEeIXBgK
Y2VqTfrsmL4xoC5xChjHfScl6E/y+tGXqn9gm6mE4S+g6pf9XTQH3zNdjM7UeJPE
EraSlUbomTW1FMu1CWhC+nwn4svkJz+O7BkSibNUDHx5H/d0Z/yU+7ya5jJYQN5X
je0fAjHtnFTm/rWSAY9uIdtrdzDdvcUSlmtzcS+9TC/mEOIZOMwb6blMklVap0n+
Yos8WYM87AKr1Okd611HwMUPeAlWDcL56uBpCDDV6ruhft4cE1q3jo6+6lzHW8H6
hTdYECGymuCEuyYVBwNbTcHlQawqAGuUIF8sChGr8ZOBCAWoUJNkcqATbW3UJdFy
qmmVsWrl2TZ+kMRA83mBhSBRRVNzIuKJ/9lHzadSzcDlMs/+kD0JILDfCx5xAZbZ
tAVOLRswq6+TpDtzm+ZdrSP31w/9Fefp4aobgsrjZDxoHT1B1LJOMrpc6G0Jfpe3
zchQrqo43pxKKgMdhivBM1d49P0gSwGhLnprW1OXp+HQrCLlCmkGao5J/ZCdcRtj
v3jeYe7dO7SCGL6tOFiJnhh2HVOhBHqW5kQ7WOYglWbFORx/bOXvBQy5FtHFBOly
Nw/kXuemt5clzoICZckUaEwkS4EJZ3DcYEOUUC09qGR3Wo8cdxQ3iB2T9f1gWnZE
3gMP2weVjcitM+p0xlmD1K3Zh6gwqNmEW9goWaxEEk1LyH2wFQpqOk54Am7ulXJJ
mc1qGjd+wWlaVS5vlt6oyFdHqKtgnYcLaDFkXr4Ihx5/gT4xKkrFR6dbpo8q++RM
Sm3rs9jPExZIV01dzKa42ohqATGdEuhxV6L3zEOFQO4NueTUiTR9o/rqPP6tIYEE
7WVKCccE4P4pKPNNuh55+KfguSxJD57J68NaiyWhqS8JUorOnQYOcRjBf0pkQB2B
GLF3Hptuuz1Tkdnn5pNHt4br+bFdfCHZ+6kDMYTpEgOhVoVJ2sM8ASTjrnscFYaX
//zDNZ4yzKt2NNrd8j+7x/kp0kJ5O/5qda+D4Xg3TUB2eW7sikjVsAVvw2g3CXju
JFoZl+fw2M3WktuiElE7tZ3s+VtUmy7wwMWkhgamt67En1K22KzU+oSN2MblUQT7
Fl2Vqc6QY/fduOkPCimPA5mFIHrZ0jLMnoChZC8I4uKWXjyC8lP+m14c/TVcj8u6
PjGqbQ/U3LCn/pb01Fqhv0N83R2j7i5fnJr75qAkwBpyTO/T7OZEjuv9nnnlT+Mh
g8/qduo8cRaRPEwetnpbiKHm88PkFu26FOGgcXUIPX/ilLyNed/ajdIisl85NPxj
ymonbTi7PedWpKU6oe9rVdoMO2xpg+MXb2p73os/rTWyqdJ6uB3GDRRYdAwxi0Bn
XvelW8yDVCKTrqHkfVwW9ng1wxTeTeboSxAkDOJDgu4m7uZsKCoR2lV0a+yN0sfx
HHJaVNFwnfqnsqdplN/WGt/poMS+6oRB0zG1qNuXfCKpUV5BrGGajrfqFyoeFBXf
mk5jdHJ24RzqRrnwi96+Vr6JvBMwwfqleaNKjhOwnj7PZSXMWbD4YEnqdGQibNmh
/CjZ7KyfLD0V+JjOX1gSlgqWYrzkwIhpXnkRtATzhCQ+KVKMkpmzOe9msdh57bt9
jOykp+0NIeKpJ7OuSU3L11FKcDexTI6Y+vZDau/3DMX/yx0aWadUX017OEMRFDRE
lytn8Hq3XKb+1Yov00mbI+TWq37AqG2hkDBHrxyIs0f8mGoUMns61nfuo2LeP5mV
l+uvKZd6VLOnuCCM0QBdrWSoAeg8QMGqMKcZ7HcqtKQro/OHVvwbJR4H2ZgAQqG/
W+oRGxprv5InGjxGTkGiN+vr+Se6R8qajPcleXDr8Kf1npgyTyy2SMa4zB9Lk4U3
zqbX1V1cG5jP1J754qqLxkDcbJwflBUOMIl7Ay75RmvDj51YqiPPVpIc6Cc1urtO
GtgRJJeZBFAirXhZ4q1QWPaV0OryI5WD80hCn725UovRAL3ksFmQ3xcIqQ0uMo/J
B0OeSQYuu1b+FAuQMKYJMPh4jub3PIVaCZYTj1kG4eLdfu6BwwD1N7tM6HKrbcMh
M5apZrMPAMG9e68DgejtxQwDqH0kg6c40H3mTxyqxGfuXsoyCS5iNJ8gBLxXqbJk
/hpgIV4jJ2VQm8q/6d1uB/usP2UrHgb10bY4jPSIe4MYdhzQTd+rIjM/h60Ju9Cq
Ym3gZdyOtlw+wArMaQIOQIC7nKcLSmCXQLY7f1Q6AO1Lww0q9qlIVFsSiiMYTbXi
HTiitinXiPyRezSwYZxqaUmfNpz/pnwrca9QEkN6qO7RgGknrVz5h3EWc6gtruRK
JqaG+n2DA3VRH4gD4eSIVI94DHQzz+fLR0GVGdQ2S+xWJuuzqlb7Gjm0wA+LZjmV
rkdw+GFSqMrMuryTjCMpb0SSnnbNDDBS1h+zgLz3cZweAurwnhD1RxqHkF0uv5DX
Wdnt6hAD4QGabMkfwQg3MPg6u8Cb2yvcGNCZT9XPSB3EnIZBbB2HXJ0Tbr5kYmdN
ilT9gmQtUl7hua8IvpfzBjbJvGYzPs7TJwATh4cDDBUCAjfZJ6H5v9XeTKcznoRe
pxQsCjxJwAaDMM9V8xOC7HYqQ6aIehCAM8E2qTuXE6l78WoePyn84P4jv0yH9wq8
/GxE2lgg4rMwzoJH9DO9PrpxEwPgPRmSjuusy6WvNMDXxXrC5aMn+Wg4Z6faJAKL
t683RU8uUEs7AMWH4U0jG0r/44d9AASjBoW9h0pncZu9xgRJG5Eswmf6EMPjI8NU
y2IdmPrxIUBDyGuZOk15zY60VqUOzbnrK2aYBg8UwfysPqGkv3nTVZ92mfGXH7PN
wc6UYybjiFq8qcxuR9+IAmy0ww65amUvWNCVb1wTjznttJrFVciqAJ6dD46r/tiI
1W+dhQ/3abEBHSN/t4FvNmsGmmOisvYvPaZyqMw+MrCOIqZ8tcOMWtlP7ukksfJ8
LLQN0jtvtdj2K7woBlry3eeGmGWpGdrHwt7cYOAt5DaMymVLRAW3jHRuJiPzB/SH
`pragma protect end_protected
