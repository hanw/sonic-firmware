��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���/���K}W��v�!��~V �qc�H_\�O<������?q *n��qƫ>�"� �hRZ�;e^[B�޶�eti����`q�<Yq"���\�I�o�Qh�0�=�}�A4	����1Y�, ,R.�z���IS������i�GG�"B<#�P0K�������z����WT�gYC�.0�� �1�B�/��٥����v/�Bf]Ip��B5��o�yk�G��h1�>b�M	�6{*�z�)�b�R��#a}8K�Zg�a�a?��c]^Ҍ�	ϫBg:�ծ��������JH<Zj����Q�w1՝q�.��_�t������ U�aQ���	2���G7��y���#_-9���Tzc\�����Hq�ټ9��oYK�P�3W�����l@|��x*��� ^`��ܺ�Z�?�]�I�U��R~τSN��%.^u��$����1crciF��L}k#�G��T-��&��I��,��۰w�~k���Ĭlqy���1��m�u �R���%���M�pk��"���R�u#0.h;y��¡����Y�#�#C������vT_��kY�<�]�sԷ3�PV,�2	d�80��+��)���7CJ����t�l��;vi��t��o�X��Nj����H�]��2�>��/
�n���I�E+Ϣ�&����IY��f�f��.!�^�N��v�m��zc�f����-�~�\���)��tzج8=��#�`��ʣ@��DT(q7���@�y;/�
����.���y"�6�GK=�_��o6� �]��M~?�/���,��D@a����!��]�T�� �3��m�����}'S�˟D��%�5�tQ��S���e��Vgse�D��Kvӗ�X�`���w�����|���S��pOA�f�A��y��Q��J��\W�uwVt��96�ԣ�o���1�QSr��o;ۃ�n/ʴN�7Z ��-I2���J���ڭ
J�A2xX5SV�*�y�2Q�xEn)�B:�����|s\�6��.��H��H���SN�;&'�(M<�*A%���V��}`-�o;�&>O����K�I&GdYb�m�^ٞb�T���˶�V��U�cIh��[7X�~
fPc��D���4$�����\�[w�g�.`�E���DN���`҅"uI]�ݞ#�}�+���w�2l���Y�9�J�2͉۝�M,Z���EL!��"
���e"��X��/?�箌^�����{�j��_��N�(%C��QoΫi9j?x��:���$�3�{��d���kIGӏ�4t,���dب&�Cz=1]��S�������y���(}�Q������8)��p,uG�5l6P=H�A+��z��]4�Q���_�$ƙ7%�rEb�wDˈ°շ3�����Ni�rP;�zmS���n�)%�2h��u�ns �K]���ۜ!t6o�!�fp�a�l���p{^x!�w�b��m�C�n�l�ɝT�L��E�R	HP�:t�ެfI��[�>�w��6��h�`šs榓6FY���֨!�6a�f6�mw�� CVP�폪���S�cgdh���X�X���D����g���,&��$*��#S��m��?����i��S|��w��X�A��VG�]p��A���	SJ�� 0�\�\�(u�j�/��iFU~0�yd�]��y���,�2��vU>Ȼ9��1�C7��|g���Ѭ��+P\}zF�|}�r�/'���� S<qxE`JO�~6< }���4Sv;X��bd���m�/�ͯ��I�)��v��X��}K8�A�N#��JR��[�<�m�YY~k���i��{�C9Y�E�C@+f�ToQ�D�������z\l�6]|�A���+��#	�arݹi	��Ï��,�:l��W�8Rռ��6�|w��b��a�鏇=��l²�` wSgr����S��c ����v��6���A��;�&QM��p��#�M�.2�!~������]u�ebz����,����{*GA��7O���๸SK����g$ɟY��7�*���B(U���[8B~RZf%h�n�3���U��Xvy�Ղ����1zsUx>��cL�
�և��!��nx�F�Vr����qq^���z1��NJ����<��z��(�o��h��19#��`��RB�G�����m��og��I�E�����\���?���i���<�`"9#M5n	onDh�lƃ���U������$����)��`p�;���u�o�{2<���=��#��"mS.��sp��A��Ң绬%\o}�o?!��>$g,V��*Ko#���c�"B���'�6V\�X��ȉ�[�an?�eF��;|�����+n�ߎ9�X�bh���g�������+/�Dviu�<Wx@e?m7��/.�},�au��Z�֚V�)����W���Ư�ƛ6>`�[�漩�^���.�)�1i�v,�O��-!*LE����4��Ы�5���z������;�����}5�LAK�?��I�mw�[�RR��jUn����H0�ȡH�7B�=��g������/��B��- �@`�s&iD֪����L�U���.�L,|���Bɸ+X'���U�eR�OǶP(�z��M[L&��p!������7��4�{"o-<�1���3�ߍ!�@�zP�v��/L�$���� |�T������mS�����X#���c����d�As�$5���J�j˕[��5V��s~���$8�����_����C� �_� };����K�����(��M�QԒ·�hOk�)��PJL�b����-��2���v�굙<	�U��F�x�?d�l�J��K�j�QR�y�̢�C�֪���@�~_�Nʓ�3#h���He^�N@yt۵k��¹+���z�1��ٛ�,�7��,��5�y#�g?M���\h��\�4�S�z~0�#�ָ�ݟ�OP��7-�����$�_<�����"u��%�"b���
��.O�H�g��=��Vp�Z��۱݋�x����srւ�ާ�4�})���@F7~�H9xk��}l�cт��6
 
����ˤj4���>|�T&p/��:Q�x;�#����!0���g��Y�W�L/U�f`�+>g��ӟ��)e�m�<�P��S��ަG� ��:؉K��}�UH4�{D�t��O�����<}!���`E�#zM7L��k��V���o&��wA��������d�.A�UI�p����`������/Q;BI��1}�2.f�����9��l�v\��J��K�!گ��-h���\��!�(9Y[�ԉ�VB��,]ΰ��� zU�����8%�$��i�4����	c0�*���RA6U�?�͵�90���sr>?��r-�1j�����`|����Y��S�AF�UH��u*RN0�1��Cqd?vT��HUh\�K�}}���9�r_�8ԗ	�8%�1������8��H��$ޑFAe��/<j�Q0NM����XԊ�*h�6��ޥ/3�\�e��-�ia�ag41i*�Hs4��Bw�[�x-�"��!QTw7��ȧ��<0���a���gO��
�p<�%k�<��k��Tk:��\�������4�g9:�B�
���I"�E�p"0#1NX-���^8 }%���=D���:[�E=��X?��:D�Z�%l�M����1�����@q��gE�����G(�Ȕ��?14�K�Ƶm#�mN,7���ՠ��`FVU�\�U�=��,�����O�W�U�(6���PS�+�Q��>����{��/�b�X���C��)�rED��ZI��)+�0���G����Mw�C��fv����{8��uI�L$ا�u��N��d��i̍{�= �N~2-sH�AO�%(�	 �Ï��^��J��p���6�?����6�����z���P�� R�`�x�c}�	M�(���R���%��?z�dD ZI�FK2�U:]�17.>>%�1&Mw���Y:dJ}'U����Pl��F=���{i6�,Hu�7�u$����@�����xU���G��L��R"x�5+g�a�#=&�IQ��,�T(Si�nd���Kt�b���H/�C�7Sj��8���x�5� �Y��)�'��|eE+���-�V@�;'�ּ|?��Qe�wϭ�V��b�x�?�5�>J^]�9#�ʉ��i6E����m�d�b����lpkd*��y_�+��,T�p4�Lwx)S��>��ƠbR�+���2�ָ���r�D�8��í�#$RS�{�Ukӻ��S��n����j��A�����O.v!?Ȱ��5U��Sz @�k_ ~M�Ε��X��G��	@Si'��,��V�h^��2F6�V?<I� �R���v��9B�&E�XG(�cߣj�r`�huHF��ע<kPϩ�t��{���ZZ��e!Ҥ>�����i��E�4���.r�~��08і��]�0#ಣ&tA�%�"����&M��[�Slt��t][�[�/�si]\����퉟(�!��K��/#Ɩ��&�,��nh�}r���N'�v ��
ͱsΌ�;`�B�:�Qtә����t�����0��)���yt𛉏��rG���N�Po
��@w�>��̫��-'!�x��<»�RSkV��k%Ԉfn¥�����\�ý���Op,\4\�w�$��N���}Ά��$S�9���a$�����x�C���z�s����b�%�eZ_��5(��8�gY^����n�1X�����P�S(�)�	��)R�)��P�
Fj-U���Ձ�������!���E(�g[�iߺ��+�U&��$���6��/��"g�{��x:\>�����Kf
�+�3{��r1�}	��$��{���I�ʺc�p�E+o��{���Xl��5�~�d/bN�~<!��r��Y&�S�SO&f1Y�e����샸�ma�Ep��縵Zб'<*cڀ�i���+�&��𲓟�P�ŉ�(d�o]�������|Pe]�� �Ѱ�����Ӽ2�{W<Q���~�ͩ�=r��]Z�Wq@#�X�/���O!��B\����1n��������&yع��}�qj8)<Kķ)�4"$I>�p�bI�iVP^��)b1�)2����%m�w�g$�Z�''J֧S���U��ӥ���>�n��X�,��bo2(�8[S�P�����+)zH�3`����#sq��;/ϧ�B�׷H��!��eG�X@�̲5R�C�ӝ�ڼ��Sv����"�\����Ǉ����\��AV�x��W�/�-*Ą.G˓b�'%!z�iW4��h"z�5ih�[�hQs�z��v`��X>�K7"�w"|r�L�}϶)�4��I�ˠ��b���Scy*��������n�+�����E3�|��̓�a�%�l� :�"PHۭP�q20��h�[������O-,�kY:V�pH��̣P�
[x�9��\�T�	�5:�f������ņ�E�e*;��(�U�D�,4$���/��j9�{�*�p��!%P���T[#��1���o�#:�0~����y����r�� �w�>l[HR4�n]�ǿ�s�'����z��&�A�x3(��Oj��S�-\i83ՙԸ\�	�)ç��>$?���G�%O�@�2yo���4GP�^�gc��;�NP�7Ve�i/ܣ~A�F��,���2�w8�Ž$I:w�4q�s:U=��7��R��Wy�	\b��TǠ�+:�lD�'qQu�P_��'��R��lE{�_*=zX�K��2v :���D�K�i���.�- {�c��=K�z��t������ڦ㯻\=�5�b�h2���6�J�B��m��2<�[h�����%�Kr�G��Z�;_v;��(˿�_�Yh�x�HbL�5���������އ���K%�hz���r�I���-7�����)%Y�7j\�a^��7�}���Σ�%���V/��4�tVW�,�De�켍D��,�L���P��#ic}Ĳ-nF�׭l������v,� �߾�Xg��-Q6��mU���»g#s�
�f���x���Xq�?�E�4�u-��"Hز�'�(��r�M_��z��S\��H|�Ӵ��d�b&ҥ�%�P �TuSt�;�hg��!�E�(�z�g����%]�gsi�}y5�n����HH�d ���}���(�k���Dj� ʾr�Nn�\k�e�ԟ(�8��Z/1wE�
�cQꖑ��TX##-��!�d��D�m�@WQ�[�����HV�8*�D�dN"@����`��>e��K��,~�)��G�W�ji>Y.�e*,���"2�������4��NT��z͐�X�LL�����׬h�9��{:8�hP���}$�$zÏ=4���H�U��d��_��W �~s��~���\ʟa_����N!G�eI���p__�H�� �i�-�<mK�����3�j�/%�$�:  pil��w�2�Y���F;��H�Q�LL��U��.�Y��
�A5m)Bj7{���W�%\��O�ۡ�=���DJ�a�����
R�����)}��F�`f��J'Gp��İ��@zp����g0>�n9*�H!k����;I�v�Bs1�jI�.�P&F"�/��#
mau�Ъ��/�F	��T�3�Y��ڐւ�+��P;����64��z:�M���lz�\���egXj:�M��L1p6QpHZ�r�5��+����O��f��R��Vw9T��@d^��4u�R�^K���h3}a����?Z��A�$jG��~P$6�1��z5w�,A�h���Ʈ[�������Vؚ�@I�q�%[bh��ffR��^r0.�i2Vnn ��;�q�M�<|P��Xz,\ktO�Ԣ!D%�<u��_y���5�?]�l+��х�i$A���t�b�O(L��i��0yC �,�.`UJ�ͬFZ	/�2�ƍEX���r�	��,�K���Zk��6o�3����u̴ U�.g��v�^y�l�Ȏt%�}׼�}V�u�-\�J̐��Ƚ�&���<�<ϊ�
��tm�H�t��k��v�̗��G��ő�RJ�*ǝxNOZy�O�?9��T.5�,��a����@�?<��H�Y���E�>e� ��r]b A���d��IT��
r{�-,�[����y�w��+԰#	���8̳�� 7�wY^��n�J��#� �u'����s�t�9����n�E�;�=��&��%��΅V�Y��ʍ�*s��U�F�i�܋��5�
6F �lLpG.��֨K��Ͽ_60���t`J�"^��
6%\��_�;,Gʣ���+e.�������P#:>���L@Q }�����M�A�Z6AF$�BG==d�'��������6M�*ꇂF�����eas3������y��%��Ԧ���D ��������\>VuB?��� �6q�9�Qbㅏ��A����=}�4�9�qU�k7gI��'�+���ܪ�����E3�M|�o�om2˚Z�y�n ��{���؄6T��Xh�A_��y�!�)<'������C�k�-�xÝ��L�]La����^�&q߄��qa�:S�$Bx�)���Z��ā�w	����JU�R(����"�_A���@�w�˩�T�@t)�dK]k�'�3-��QAq2D8:nuۖ@�?Ǝ�̈noyg�aD�o�W<r�@��bɣ�ʹ���*=g��VT#���Z,?9J����&�A�w�����.N��� �J��A�����U���]:�Y&Έ����L����1�G�$�����v��-V�j� ��N�Q�?�o	�����H⥎�͗��(��S?=}A�Նp����
_�6Ƈ׼8��j�E�rM��K�D�Zۗ��͕!s�F���i�q��'��掋s�E�%|.�ќXe�x�1�x!��9����9t��1ۑ�T�E&��DPe���]�ŊC�p�Ϛ��q�#�L���z��u��f`qVT`��M���H7�H�Ӥ�I�Ŗ9��%���{%7vu�}�����A��YZl��1��YG�@��'��߲z������f*L�0��7�s[^&��t�bc�R��Ռ(�A
�����՟��1+�z��m��d��ʢ��תn&���F��u��DÂEfs�+�p%8$���ρ'�d��a�p�`�l�V�s��}�KM���H�V����K
b����<ǯ�A���x�LjC�e�b}�*��ktYC�w��8�n�H~y����u?���m�d��b5h)H�Ȳ*+46�ǒ8���!�����1��PYPY�ǒg҂ /^pϽ��N.~~��\���^4�xaY�H����<�����&���5����~tl�og���=�i4��*T�w����Ā!ѡ�Tj��O�7��?���kv2P��(�ǧId����ί�.��e�9�1)��k�J]X+0~�l�4��2� �ϳ�)�����7�%��~�}��b�Ymٰ��@6��'�ma�j�:��i9Ұh�x<��8���'���fF����q4#mT�|���5Y����oӴ���wL��g:
��3������%ʽzJ�_S~�O�l���U��v��fX=J�9O ~��+�2�+&x �[��Sm�>�����w�<�9���g�7Ls���,�PJ�y��-K�?���Cr�Ќ�C�l����7�V�j<��v;!ڕ`דҜ�kg^��V�J,����Xb�vVKЯn�g�v��&�f����H��B'���5)�R�t��QG~u��ץb��@>��l���H3:k'���D����~�J�t8�[0��˗p=���{�ѯ��)8�W&kj0T	y�k�:��}��m�����.2��a�Pr/���{n"����ǅcH�"ɻ��h�O7�r�1���L����;���<.[EA��Ps�>�Q���ǁ;���i���T��B����T�[){��^s�����	��Y_�LA�<�CW�)���-��~��3��Q �N35�(�Ӈ��R�mH⥦�C7K�I"6�A�����X!�a�b@o�M��ߴ����(H�yE�k�S�!�q��a
��Q��� �ї������bh�b¬K>��TEi�u����*�?�Z4�,֠���e�<�<ޞ2;ځ�0�Ѿ4��gM��4@ \�צu��GF[Ly�R���l��(.�ε`UtK)B����B� �ܕ^!1 Ǉ���\�����mH*61���3�s�n]��=3�2^4��������a�[A�s�&X������Is����������ɂ+~��a�(辩+`��1-�	R����#u��D��SmŴ�)�C�X�lUl������Ǘ��ҫ��.�ç�~�7}(����eo�"���>�5T��2eD���푶�R�3"�2;��s(0�=�J"���ʘt����v}�d�[�!���}���A�]P��9^8��݀�?����ׂ���o1�g��1�m@_�OJ�p� g߰~i+�s�1"��g�5��H�7;�ށc�E?�_��w������ÈW ���:��a
9}�︶6�eE��v6e$�I#��1#�y'����HLz�ǝZ�2�w��0�Ljp��UN8�T�[W��>.��j'����ߜɶ����ң*Youm�21�׎��HU�0��?;ϟY��y�S�qP�J�MJ� Ѡ��L ���#[��a7���D��`�7^�g�S8-:��,��9�@�f��=1�J�L�7��$Z[��o���9��-�iV�f)뻶���<�2q˂�6�E�+;5b1A?�v���L;ʾ��4'��� �sA��zf�.��XZ_�N�A���[Z��1͔Ɛ>�SL���`C0oƓ�	�`���\:��x�9ޥ��^u�/(�Ei���W�G9cSC���`��@F�����^S �a�����v�U+�|���g&$�x{��G �c���9B
C���|v��5��X�X�ُZ����u�v[���+`L�n�U˹�,��p���?�X��>��/g �_W>8���p	q�H�=�X�ŕ�3�U��
�����3��4̓M1�OH���g+�L2�g(AR:��G�G��p?��|�9�������#-���z��r����K�y��|꿴�M:C�~O)�j�Q������(b,��	L�ݯ�۳"���}�N&X�=���!�w���-�h"��}G+�7��
�Cb2{����t���}:��Ӭ:OM�|�eEr�w�UV�2�l/?��0\�u�E(E� D�]�t�rC�؉u�Œ'�[�������LL�~�-:��<r��6�:%̐,�zr�R����h����S0�f�n%X���,�!@�����,'6���^��csЋ�*��])Ѿ3=��@G���az'�������br�����E��Eή�,�MdX��ʗ.�}I+n�)@6Y��-x�e��Ft��낾\�اa�mo���#���_aP�-��L�.�g��c����cӛV����%u�]��,;�H~�uF�69^������F�<[��_Np� ��
�!��:��؜H9VN#�����8�����������Q@�Ի[����S�.��;���jڞ<˹�&Z��#�/%D;x�%xwY�쀏U�|�*�Y���q'�3�q.�-��/�+t�Zo$�4S(�'i�U���#�[c߽ $XX�^V�}���Z����0G���+#��e���#h8#6�E���Bf�iZ�M�K�	ƪ�E�N��~M�O�jk�׷��}�4��R�����F����]-m�H�oaκvJn����G�Ue��8�b�V\�8���8m �-RX%w������mz�
0���<�$t��<����CCύ`@��Wy���OR��-Չ@��Y6Kl>oZF{����q�]*C�ֵ[:����<0=���h��<v7@��|F"�+�����u'���韁���!d���[�YΒ�Y�ͅ�ғ�g!���EY��A��΄�2c=�:v����>��X�(k0�
������q�
�x�e��>�Üd}�H?��e^'�G��c��2�t~BN���A�x+�	�{����<���rv�1�q'���4�5Z��W�3{�)p i0��m�V���Ţz����f5I9��q�Ų��P��R�1�7T;����X�*�l+��(�����5?�J�!�r<{�c�Sx�x6��	vf��"vH����v:wLc�������n+c.�r�`�I��rX+G�f`J|�� ����g�p��[�L�� �7��T�x���Я��J��9%���"/��m�3g�豛�ϼ���Ø`�����[әI��jQ6�����pX/ve㊩tځ�z���U�8#XO77�m'cR��ئ��E��%7�?I���gx�GL�*X��K�.�;2�;şQAɇS$��3�����aS#�v��{��~���({��Pι��l��L����i*<��e��tqy��On�v � � ��-Ȧ��i�?��q�`��G�� ������<9�,Nk�ȼs�I�-[�	1�K�^{t��'�1�co){�)c��8@f���´8����A]��\ �/��]�����kT��{h{��~��DTYs���!�18�lGi���5uՈrM�m����R��5 ѣS�wM�wB��h!C9��.���Z>^F���&[e0�F�:�y��r���;X{�[f���_3U�*��:�n���|��ম`��{%�'�4��W��E[Rfp��q٪�/�� ���ղi���Z�ۼ;�c��	c�(z#cϺl����9ɍ�}���3���`$��%1d��}�}�-��nó��Tɞ3k%�oE���=w?���m��R33����V�Vͮ�ٸ'��ӷF�>M�����{"9�.�Y���P*%=_<�>�W2a-cǘ�S�s�F�[AWQ�r���?,6�m_�Ц�}&O�s(�Oܣ"!����z���@]M*��	�6CJ�9��Bih���nq��s�'Bts`q�����f���2�p�w��T�OX��&�0��'���o��>RD�pl�z`��D�{� ��4���7�1 ��n��Bj7?H�����*�_��nt�S�1�{��_P'�
|�˚��_��n��0���L�F���;z��IĴm�]$��<��b�~���i-������`�˽�I`� _���|�V�^�ߡ�v�>zH6yM��I]��8�0'UX��d��W�>NEv�SҕS�kq3U�_6�ĸ[k|Z,�Z7��;zܳr�1��NA�>Q�L�Q��l}�w6U����� ��KՍ��kv.��߉��Ʌ�����}m���hփ\��_��6iVc!�qo@mv�q��U�8v����r��æ+���\S:]q���xчP��Tt�j��h��f*����nN4_��}��&^����Ɔ�/,�)�5�x^�r5��a�6��;���wٔw�h��K�)��.Sޭ����J���h�`����#�bK�}q��<C��v�p�_���kJ��`}�Qg�>�Z���ahW]U4�LV8u�D�(������ ���Y���"�Sv�Q�V
�#�)�
�O���JH�c��<rm(W	в��F<�P��I:/��`t��9tdn����L�ĝr}�,_O���Ŋ���=N�w 3EIl��b���B�x͘� �ѐ��Y��>��#b�Âl�.E6��Y�%zE�@Æ�0��>`8P�̵��F!�Є�&͊��R²���De����ci��u>L�ܤO�i�θN`�"����V��Q�1��ُ���`�tw�;��&���7F��t�j�1�s���W��^UR�,\�� [�
F��}c�ӗs�b�.��Zp�U V��-�֥��O��~V�B'��׫:Eq�Va"8�2�T�?�ڼJ�a�r�\{Zp(D��3�V�Kd eЅS��3G���^��Qp����н- �*?�ᨫR����ipe��HNl��i�uށ�8�\��p�i�e/���;�2k(h�x��hт
�����2�8OY�#6��)(e�U�f�z��&j��/�����k�5���>����r0v�}�&����`V�*��*땚��$�Q�삾��U��^/=�T�%�q(���Qǩ��
gO��H c��<�
��	~�Y�� /�w������YC���?��k<�_��}�K�\#����;)N�K�"��4/������`*�&;��k�W.�	��,���uN����9���&@�� FQb��r\�6� ��r�u�h$��̓�x^bX��!f��oD�b �8��rq-xy��K�*Sa�Y�y��	A��෍!��}|U��8�+�)�!�D������ܬHOw�j2�
e��hTf����8V��h^R<�%��pxyy@M�0�^5^qk�H�k̬x�vQ�Qʦ�@J%|��4��e��`�f�	���,�����#b���-�"�t7�R�ײP/E�sX��PCȭt�t !¼�M&O��.�y�h�G��$5��j�9Z`(��΀�>�F��Rљ���z����?U�x+��Ǥ��|�4b��{=4±F�?=��3��XB��M;��8]K�J$����A��%ı���!���x�)�����Z��/f�$��V�0�ɧ� c�VT�de�;�p̄��0_���5�u� �]`�
��b.�;(9���Z���mp�C�l�o'�!�v�*mIw����v;��f#�^���\k���|�C��7�;_]@�q��������G��W��,��h��/�k�D �c�'�"+��q��+Z]�r���e���Ą��$r�T��{�.�:�I�
��#�r�^Z[�tӟA�2������W�=m��š���,�Y~��R�v�d�����U�NL#�?�6K����3��H��Y��sZDm$���d
�����Q�S�@��0b� j�ni <HW�LY'�A㨓ɟ�Ûpб�F�����| ��J���m�V�o1Wv]s��S��`= �BlE��!����z�q�B����K�&�f4�4<5LhE��bt�L�hUV��� Q�0����PG�!�gD9[�Qw\��I� �c%�Pm@��s���8a�Y��)�/��<T^kB;]^���-q���Dד�������lpX$��3����С�r8�	�k�rϯ>����N�uɮE���ɫ0�S��s+�yS��-��6���d'��� H�Ȕ>��us��"��p������ډ�R�ko��+	d�yz�9�7��]nkBL�} 9+�f��UCC*���}�/Wo+O� �A��UY�+m@����(�:�T�QE��@x�S�[�D^�D�^jz��ㆺH"#| ��X8�-y�3������lIV\NFA��&NP�0Ƈ�o1���s��	B]���tG*_^����<_��	w=�_t����	��G��>�YjQ�e�Ô(;glKr�D�]o�R��NZ.Y:R:U�Ts-*�֪:��&�A���`f7�Ky	ȠpMRr�=�T�<��=^��P	Z�Z��Լ�<J�@6�z��5Sq}�0N{�	��r��3�o_�"quv��`x��Ƒo� ��D�|Ģ�'ׯ���y��k�`����m�����6��^,НI�c�#�ݣ�ݣ��#�mi��o�&',���E����8�m�/\�| ��1���<�>�ښ���T(������9�6��6@�-d�]<���2O��3�?�S3&O�/:����TB�s.���R`���̆����A�̈�G�x��WKf�fNZ�E��צb4�H�q�ء��|I��x�W%���V�~����*1M���FL��|E9�4p�͈ ^�;a@q�3�(�܅~`�J�?�T�R,�N����� >c=��;�JoַfTU�������bhvj ޠ�;V�����R�V�m�p�N������k�Cn*3��l��`�7�biSc/�C!�`f�/�@�+c2+}W���qE6����z>}���4�h����r^���A35;ΐ�n��&{�g4��*�I�`�S^"�eaO��duR���f>��N�?��U�[���[�{5���+����^U]�d�T��2��ܮ�n�h�2	˓�5� ���ոW=���wց����_�J��Bl7c�sb�MY�ZJ+Ζ)G��Ք�(��������ȉ�<�y>�J��Z������?8�'����C���_�b2o��ȯE�Ih@�� �cF��7|����!���Y���F�D1��˕y��1V�ԏ���P�YT�}�]���+\2I��
�������E�>>����~+1-s�#�8 d��\�w�6RԮ�Pp�zx��eٱ�C��C���]����R\gy�����4O����45�VK�R����M-5�7�V.���.u~��x&���'�;~П# ���.�_ K);��am���
O3�<?�q�ƽ�|�ꤴ7&m�
��YCY�Ή�d�r��B6��g%�Ͽ;���G�5ᕔSÈӳ�G
���G�3�)hP�?����nj����Ĕ)(��~g�������u����H�P���xy�2�;ڨbr��4�R.����9����F�O��V�h	����)�d�iUcZ�� ��]Q��)�gkBi�N��8h��9q2@fv���k����d�*:E�G^�!���v�=��I�rD"Vk��}�L9��F�)�#�iK�N
`�0��q�`�䚈���@�
ad�<��lպ3�1�Ԗ ����QX�m1�Ε�`C�r�驠�K0�U~�\HY)�H)��DP��<@U��U\.�m)����_�`Pr�<����H(<-j������%n@b��6DY�e�Yp�58���k ���g$8��v/T �UC�݊���~V8�{��s!!�P�ﳯ9�2���K�g/ő6h�%Ҋ��TR�d��S�4��H���!G��g�����ƀU�MR�c� Z1����J�w[�ҖS7u��1�s,�^j~�b6gs�~���iAgw�eΙ|��=�Վ��-�4z�Cޑ�"!��6�,f�'�F/U>$#:4Fq`ݦ�뙥p�0�|�(�(q#RQRj*����"%���a��7'�bw�OHw��"$Ay
�+{��MdQ�G3Ǐ�6���� 
j��_�=���n�3q���	P}�����!ɇ���R�x��x�!_� �Bbj�6ʷ���~��T>���B[w`a��i�e���Yxy��O8mƝ��_���0�J�g���� K����%g�>�ZVH#$/�I�A1wT�X���m�ի��b�k�	�J���/�i������������yLW{h�
�صZ`�dV�Vzuy*G���^vL��ޤ-��g�qCE4m�����Ꟈ�2�Q�b��0��S�~�u�8]�����_f��L��J%��ܺSy���(��M���`^�`�崦��5[>�u��	ˎ�e��6U�2E�b�ٱ=У�:���w�c�n�R���=�r���Dր��Pn�>�6�b$�H�tO�k�}v�� ��e���q-��
 ����Ū$��8�4�[󫤧���]V���G`������������(��U�~*�5W1�Կ���Z�3$F��֊%8y�����z���������9b �ħx=��R)��5�r����c}&�nW�/�$�Ӈ>����(�Bl���Ь}�B\��n�sH:F*�SE=;}���9@�Mk֫�}$���09C���&�Pc�Ɗ�2S�B�����p��n�����ڗƏf�p�"�սi�E�e��gw>����%'N�O �i�֮a��>�G�ߊ��w�\���;d=>!F����qt!"CCS�*j���s�荮���Fp���#)�����+T���F6y;'g��Pn�9�x�bȯs�?4n�{ 2�)o��W(��n��	yhiFz갅<����d�E��[RP�3!����\�T `U�+ó�Ϫ�h��a��X��\c ،[����{''�Ju�P4���7V�u>������>u�;9���c�XY��GF����b$%&N&���wR��r,����6|�����[�o�O#���9�a�A�A1�8_�H?��>Fo�����#�Ib�G}d�3	$�ˤEB��X朅}
ާ�dQ�qv�e��� ����,��I1q��߿f�v!%�l�L����ű/�f.�<����/u��i���F+���y�U<�kWE�	�l���������I>��q�S��]���5V�Y���v���6��	�SeGI�Do��e&"4�s�@�è��e�߹vB��q��	�����\��g6y�)7�y-<�a6��=⤷�IӠ�1"���K>�j)r�5�ĝA�ݍ0])e`1%�P���i����I;7LW� !������$�h,�+�� :�C;�Ɍ��8*�*�iBD�	���=Z4oNBۂ���R����� �ǖ������/�7w�ϡ��A{���,?���u�FR�㪡M?���1r?��rmp���/�i�+��|q�2^�ɏh��Q�w�����냓��7�v�J�����D���d�$��m�:�!��94|�G!R�m'�55��ӑ2�yӶP��#���H�e����8�y��$�)�m�����|66$>)�F���)D��Y��-��!�������t���Лd#��!u��;�[�fA�o���򊷞����Ii�`�*t���W����`j���(˝������6�\�XMOU�(#���&��.�l�Pv�ѻ�i���
��� �r�k��1�<��pY� _�2�>0���hE٭ȫ��)q��1>C$�,����>V(��L�uh���n��Pf��#�;�d��i��S
�}���mù�;�A��1���&۪���|����1�j �p�N�~B�<P�<�#c1�^�ﺂ�������^ԥ��f��˻K�LE�\���sF�j�e��M�,����v���<W�X�DR�-@SD�7G /@N�G�W��o��9vB��Bv��,�lZal�{�Fݽr)��4�z��UJ�bk��cd~ut�wc�Ii��ڰaSjļTO:�{A���s9"��z�5��q��u�9�����0�Q�xl}�_�Mx\R�U������G4Q���� ���ʡ34v%�<�	K��s�B�� �G�ǯ���7~���N�p9"��;^iz�i�KHUK�S����<��9�
��iO���sG]qg�c}��S��g`n%�K��ğ��`��S[ ��[NP�o�xq+�(���,�<5JU�H0طUă��>�׭g����碩wJ�V��x�;�V�*�	�v�F�)��i��z�b��Ӟě�����+��Fd�qVp�÷Q͆�R'��!�E���L�7V�W�2;�癝W�Г��,/M.�i��v��V���q��b�<8$|����I��941�~uzM6y�����^�6��JX,A�`Y9*7K� ��a�7S��ߊYS]X�5�������&Ym���_��TD�sbA�������EEr\�{i�΄���&� R? w.Ƞ�FG낆n[$�u���z4���!,�s��]c��u�����m��.Q�[��W�7b��Z�wX\#C�6Ʉ��a�o�F6����	��o=�7�)z�`S8�	��"/@�z���tb���60�0��^�ʚѰ{1�,���e[�usm�����H���g?[�]g��aC�?�zvn�u��S(��9S
��%�,�M���o%A�'@T��}��	�FOrW���J���CA���1��\�AL���^ٱ]�`)i�Wb��A�Y��̲��A���(��I;s��}��h���u��7ҿk*��JZ\��4t�{f�$OϦW�!|%�&VI}�7�W�P����nM��s�K�P�/Ro��
5u�a���E#wDP�g��c7�5T�@���̽�v�U�4��θ�7�-~���� Hxo܍i����I�.^�R�'���G�����q����}51�
��^�����'2^��\Ct�f��7�{�%�[�B�Un�l�@j� �F&�d���!���7��
#����+n�V�{��6�gUB���`m[�9ag����4�Ӌ��7M->$CH���"�ĶKI6��J68ŠhD�k�9�'0�A7l�p9#"^>�����)X��X�Ms ��F�s���c7K�1G�Κ�5���8�a�E��!��x��&��f�D����Z�&%�2��H+����epVp�"M��28d��kb�����x2+"�������u#��٠�2�b��IU�������x���چZ��T}D$6�k�K�Dt�(��˻�D�a�bX��+u�� ֳ�ȸq���=�b�Q�뀣�q���V�����	�'`!�$CX2`jU��>�h|����:������*��oJ6�A��zܣ�Oϕ� ��%+K��X����Z!%^i�Q*sk�n�e��������� 
&��?Dw�d=/�NS�r�[/3�B� �Q��9����!a�)Uf�Ifx4��Z���qx��+�>��{�.�F��o.@jͰ<�����>&�j�s!���1�a��|�8�r��X�*�<n6M���.Z���lZ��Vt;�f��
Do�Zp�Z�,�/ڵ���vy8�㲈���g5ޤ�Y|�Z�^~�c*�������썀���25)�����[�@�PB����۷)�����+LIp%���m[�;߰NQ�i1�qf�v����}O=���e�ׄ=�(a�K%�A @��W�7йP�[�N���꣄��h�3DE<>�^��}W2,�[�G���玅�]��r �"���"l��S�t��8Y��t�����,VϺ'M����:�@W[������:�g�#��}_���+��叚�R�k�.8�~��2�Ǥ��G�j׸�!�ϐT(Y�?%wT:�����?7��v��8����S�j0��Oq.��7���{��(�����1���ʞ����$��#��Z /�C�lN6>���sf����Cj�K�Ի��RĄ_}��L-,rY�bW@O��ܴ���^�G ���5���n��xw��"j��=������Q\\v%� @0v4�t�Ĉ��$�C(��%sB�B�Ȟ�a��_�� �<_��I�\�y�3���p~��c������t����o�l�5	V͞Ζ<�+�'c�1��G���]C���h?�r�/=GP}�+����`}�^z2 ���3Ii5�����U�(}�}#��G�w��'�[F��|�yK����H���"���m�GD�_�VT	�Xzۈ�5�͆��m�ΔZ~@
X#V�&�C���c�����Y?�o���'�M a����O��_!&����o���:��OE8�d��c�Dⷖ��19���vv
4��v|��^�����k�eUM�#�Ka�vCɏMGw����[��9��&���u���3[�* W��=����7&�b��(D�P�":�0'"JC�iG~��� ��Ӌ
js"�zRև�B�+<�����Q�LM-#3J���|�K��c�~i��&���� ��t5M�jK������wXv�EiR=R�Y�l:]c��K�Cކ�.d��4	f�9 �[��/�-�9�A�O���`Y��@5����]�5^\i�U�lI�*�w���Ŷ�_���}��%⾐�>�=lL�Ie����ығ��K0����.�(y%	u�>����ܳ��A��ċ���/�Q@-�>7�lY\�?�Tzy`Y�19)���.F�@wcg炥�w	+$�	�����x���Y��:9�lbdv_��B ��p]�u���앯i<��t����Ӄ.WC2VV�A�
Ӵ�s�N]�ޖe'�FV�`8�O���eM�:w9pi�<�mL��͈�+��XEjjT A,��6Ěo�S��LŞ�t,�,w��_pܮB�%����a6�2�G0ȷJ�}c��Z��ԁ�>y��\�U,C�/�0&��`g�եV{����~Z�Iޟz��S��m���r��
aH\�w'����54��$��F@�=��O���ZK�g�FRn�)�*��9�~��y�&�j�������~�u.��9)��~�; F���-����M�������S�k'b����]QO���f�q���i�c��&��*���׈��G*x�G�]偰� ���2-C�J�s�/�V�,�P�}u�҆R3��ۛ;�+�u*��50p�/Q�����vGAଃ�[�R3��̽��1�Mw6�������"�m��Ca���=՜����,��1Ca����>=+  7f�G�7�&4�'���&|g�����HX �f^������T��	b
SɈ�ԃπ
ڐa�KV�Q,���7�\Qk_|ҷ%[�VCd`�g�U�D���5�R��p���\���~�Q����LUZ�BG�ɏ+yȔ�S��L����a&tFv���fKKu�EC�#ٻ<��H#���Tv|�x��E����I��ӲK�)�����!�|�H@;��^�%h*re�Ή��s�0t���t��>qJŲί9"��S�����O.�׈���$�h)��_}�
���/\%8�Q62&ް��)Ϻ:}T]H��Da%�t��9x^�6��� �g���"�1�sv��C;A��'Df����.�&Kډ'�%Z�JD�EN�h䝓Hߟ���36n��$�d��e!3�Y~B����h6/�;o�3sY
��V� ��0�كp��R�c:pR�a�M�w��h�?ڐ�Ǡw�|�¢<⏌�ë��x|Y�E�%�D�6�<)�M�~���Q��ov�\@�#����MP:Ƙ�p�pS�o�o>_�