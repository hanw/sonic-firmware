// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sQTqdpD+2CKqExMuEQQACvXrm41ibygvIDCzz8kTdYo+einmbeo7tQHhTXZDJfWI
tCK6/yFiXVQNTs8unuc7nmTRa/GzgwV50sGWr47w2zWlinSW4uUquwGZ6KBjd4nG
a70psZkcClRw8i9pe4aRqsSqG12670cSrAjzopOV6SA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2496)
uE+pNVyrFlfni1AvlY9kR4XxRGfUpmTm7yAcov5hJ1PlU2d/R1walFws0NGzVaEB
7hijgq5/ITsee/3BjAz0MnEhyE4X7dq4N8NnBFMf/k3tGGGptIQQWdRPhlFRHzgc
15jnwyD+/dfIa3tGlCOJAJbuJrv5mq0XJhPhQNnJDixpTMU+74GcQG7Cxkp2RqNQ
B/TRvLVcdQel76pkbfIWDX7Co0pV0mErCB3SgksMQS2x3sQXoLHgngFZ7lVN7CN8
MDmQ9ImSlJqpgOk+BZDRvOfU7GTWawYMusJO5IwWQZgeMFG7x1rYbcE8fLPksXnQ
AtavrMcMcnJGcCR+s6wirrUMHZcUCcsXr8W/KYJxKrWT1mVsn3/lLAgu/FLgOi6y
bjrpDgu6UC0jkkFt+8ufgn3HfX07iNN4vwG0JB+Gfk60XQ2MXWf0nrvNnPFVm9m1
uqd5IyyHJBZoHjWY6SWN4SJ4RDxkVMHqpOX9cDwlVErlF1yGLlzGYwubxR7RWbA4
ttZr6WSVxUVi34n8SlsZxwfncNvw7Rz+jP7rkgHFH7FahtfFnvDYalG/zqhMwfzI
HvHQrvTMneiVe4wriuFkZCzAj2dFtMwRX06m0xhwJFUT3vJawq7dklXOY7tWLfh8
uQuK6PfgcM34x3LAvWtNLw5NImRlhxITiUwUNshKZn2Lz43kRUAezULE7FYNUSBi
RmoXHkpcK/kE2yOU0aUog0BfmgUyPxhDT/weQY/nAap3GChVeVSUUvowQZ3t6MJS
zKjcYHsuUNFkDhoXKSF1TvI5kRhYbaX16TwfCBD4PQrFfnn/KYF6D1YKvxNNO8s8
Ch+PjjeFTpYJvQIKyARqIg5UhHCsV2H6w0hPt890dcAS6TcEsOzi0yytnRuCdgyr
CISpl0M7/6sQoowgy7QgBWsUmCHfz7+Hsf9afrmWueGLOKgP2N1s2B9dYum04KNU
7OPGuOzgU7EX+qCJFcT3nDeWFhZEMFhNOHVwNWa/AFZKo7eiMEk0zVbqAIbReEwW
J9uhaGmOz2pupq0yxB4dGn2GS2u1DBEXA6W2BTOO2wogGkR3VOOus+ubXTBnZteM
9RhzEiMr6GgyJuVarfLaqGpA9CzP90DRHVn1lPeMDpp7+L5ad4Or824UFE1STjLF
CzaUE7rQBGyumUTfN0srEU7g0tSaKfYKczGlgVSQ0QQJZKcAViCB1Q0zdbDb6vy2
9RL3S3ofTvhbEgzUr2TBcZgD5bs2UgPUOgRKBHkLDoTYtZjT5aEIXaJlOQCz0QKQ
ONM773okL3Wz+xfpKE7pIAJx3ni5W1VmVwWhrAeI2Fmv9hGn7pG60c5xh7SZ/g4n
67J7nEfiEBW1zuvALw0saWdpvs+Ser5A1rU3cfUUhucyCR8fKWVAmHRZRBlh+947
Myh+/jtyJPD3An4TWoicfvgmDIrdjJzvsXQUk1jBqgA6/avrtb9H7aLZZoxCneUc
p++AhvdWsFVioPgY+2lseSYx564OR6biQf4p/At4I2z5Sed9QlnQCTqRf74qe2pE
/djh9SktolkQze1cgh8NSg4BgnUdIayciE59Re4ObWOcQG1dcpJCWl1+wczGaBsq
VPWqWxzR5YzW6Ba505x8LH5lKPiZikLcyrdM16hTE1zwX/c9fKa2Br4zlLf2pFjA
eKxIRXKPm89p7nhJr/NH3NO/rr2BMMg0vcsVRUrfnMEvA0Ylj3Ymy/lcF71imWry
3aJ6o9eEUX0Vyv64aqcRj9WCITi0mZBLJf8IY/0cNcCTyqi8znjhQ9O73aVZ/Ltv
GC0SbvcyBH23WFW7eWrUsLuz6yTh0hHZ4C9o4DZEXi1lBXcPYCXPJi0E1Lt4D5Sy
l1BcrmbIOXwyXlvWI3fSn7jTp4I/0bjk4fcJwrsB2RVSldxmGaXu2kXQIv5ge7oj
ZKLu4pivOLkjc2JRAINBgXrXTARMeA98yI6New6HdVRJCjRGRTwi/UQK+qQzGOGX
5yTY4r0i3g0O02iwgXaSNBGcABR0tK7KerG9lyMe47oqSYIsghMtGW5OdhAprD3C
Tt0iZchrALlT2hvMfcnnPKdLr8nv8E69/opvkNPo4WLKorsWE8KI0JvwjGVRUbTl
IJiGGjpTLXj7aQHf6bJpfkDRgClbUpdFSWEyQSM2JAJqfL/OHyTUr1b4LoWyZujZ
tNCmujqLhCGJXMgvW45KhaFBupHc2lV6RAci/CdmZBlNWWoslCDnBNoHmeTPpesg
pe6P5Zl0ynEwswrzWLc+e3SdaVeG1f/lY4zcSnpeb1/JLt4EzV+71o3nY2tG/L5I
TE02UXHUiEpq2736m8ogIfxDZ4Jx0ZY+Fxc2O3dUrXVJWx+6I0DTyKmn34Eljqpu
F9+T+PXWDmsdfRrtr0p2ywWux9kuD6zLemIAmII8mBLptgSXvQxNFVFqmpXyvy7x
eT0HyfULQHUoJ9J7yr+aBpqp7RiIDG57RW1labDJoPRqULPtZrZKCzlWVlyivIy0
6k47LePor/I/z2XY2dYN7pspl0eia16ta/kudFFoPtgd825sn0uqpSW57MusZFfi
dA1SF2pXyTOVl8eawfLqKjPJBVvHpkMYkDSK94ejq7eChJ0AW0yj38fAr6wIMfeT
4um/+sYYqP2ivDRJGBMGvu5KPJVBLABugBBuQ0FratjmV8OzxHbQqoMX/s/g3paE
JvFYwEqDDxK9BmTsy5hHQLVnv1xIonoZqZfrvMtIX4tqkgsrs+kaks8xqxp4yrHJ
ET/Mdn8KbUvFUnSlC4qY9Dw7NPUfat4DReoDvyeDOXrapGIjCGDeubdrrg0bRVlp
P68fIM527Dj67KP6KMnaEg4aP6Utbqltvkl0CLkVTv1HqdB5TMg+UyvZwAVLgWev
EqokkPZFy8DbMpZigauAovV1vIOpU1Zw1uCya3OA5wRYFyeSpkSJxQBW/4Zv6MpV
wCc0Q0cBNpJA9mKY7J/i4uqM5QFBmFJ/CDMObrXLgbZniABxhuPTvSar7tZrR7WX
Xb1cMayBNIqx9jwGDdUEBFQElScufVlm5RcFM5ZbjnIEIuZRCfMv7YGpxVAjb1p4
JgCp1rWpahStTvG5VA7L7RuGaWHSBGc7r5BDM0+8HBED+qE2EyByK+dI2Y+BPmQt
n/pxzg5JzulSo+pFJRSD1BOb7iJMD488XtNDeKYiLlJdrnNSVKC9eYFDZzjl3Py6
1nIMMsLcrkY9SvvUJMl7kS71DoBqP6eIVrXb0Va+FHteNvlE+pYsyx6V1EpTq+pJ
af8pZSY58LgN+NcNcaT71YbvOesk8lHjZer/YdcVN7bRA8kcHwXfXVA6neGJcNJG
`pragma protect end_protected
