��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z�Y�$�Fe7����m��3S�	R��f��&�	�F(�RZ�� F�9>����E��4�zi�G��{�Z,���WI&l���(���5G��1�kR�c���7H�̇�.dfHI�#��Z��x,�����c���#�ţ�\A ���%���*u�:����o�9EHN�PQ-?�3)��\����bYŮ�>g̀�H��FE��KQ���L��v\w���R�4�_��!���v�0\ׁ2�TL��T"�:m��V�J���e�n"���%sn�Ep?a�G�L�=^d`�^�dq6�_���!���8�$�լzP�7s�;M`+�[�=��i~�`�2������(�y8��c�A����(�<H�p�`�KW��xwI]����q�uSW� ���$!�R��[��x��9q�!�y���Y�[N-Y��T��5^	���3�.0�.E4s\�I��B�x�J��ۯA��?-T+&�䈠����"ᾂ�z:�H�?usy��m%�/wL�M�z��:s�����ݚ%��)I�v�8e�9���� �G7&���� �'@�

e�����7`
�v��s�P`"+�%��0�k�&ٯ:$���G������rr�=zeS�U�k5ٽʑ�)���	ѻ�D���h�������v�~bW����=
��"t�t�]jo��%[|�L�V����e1�EN��U���k0��r2.�f�̡�Q񈡯�
R�1eZL��-�5ki��?��g��q5/�;��������o,���e�7L�1�8�1?��z/��(��
��Q��n_k�IHB��ʇ�k���z��P�(�c5a�$e �I�/V��r3{����w�4�`�;�ݔ�֠'.8�y_�0L��W��x�\�abt�P��b�#aW����e,���a��#gZkh�B�i��dG�}Q��5Ϙo���_�*��^��(Y��˿p�e�T-B?�bO�U��E�8:��R�TTL���F?�2��#�FF���a����؞Dm�>�xg��OG��ذ�����+��w�3�'���&V��Hh<[d�e�ZZ�qX��8�@�Ϛ������s����v��8��W����������1%���4��sqىF��I�^��f��!~$>�qzc����:��(m��t���|A�n�Xk����n���s���R�P� �����.�9h �qr@�^ޯm��0N��A�@�e܏�>D�A���
7���f�(���[|���t�LN-�c���-����^����f���볤�m����hv����) ���|�]k��I�v�K�3�PU�{��9�N|܋N�,�E��)�- :�-�#{�ń��r���M��r+����)g}��PO-x@�,c���N/J��,w��n����� �[�Z�0g��>���ՃV1[L�p`���p��c��n���{u��򨈾 ��S���t?�8?�" #�}��Ep`�ti�I�Y�B�q�{�k��uj>���2�aڑ]��u�uQ(�~;de㺊���ϋa���H7=��|�U��)��q�)뉞��w�$��,k�e�`)y�-�, �E@���"kx���?��%�ʰ��|��L�6�0���o���>Ln�g:��dq���\ǫ��p5��-��h������K�)�� �*�Q�j��nl����:Q�k���n�Ѿ�x~�,��7O"f��/zk�&M���2��)C$r��aN��G���
�s�惝u�I������)�6�`����1R`}"�J����,t�����s�P�
��E	���M�Þ��і��bZ�uNyп�:�1otEr�Ĩf��8`�폩P�E���1��-Z���,�<A��b��綄�$!�u��]�LZ�	o��P���0�VV�fUS���g�vۗ���>�w��z�.S�Ȭf��%�����Z��wŤ�����P5��ˮ��G��7�t��yG�v��n�\y	����%E<-wY,�z�Ƅ�ăd�3i/#8&4�h�}��-=t��n%].�R6����:�Ո,�>y���p�5�V���.�6ȍ�V���ǚ�:�K57W�Nj�����}��7H,|ڦ��|Y��|�������ZK����:U{Ob��(>�j�'Ę�S��]$�.��I�>	��v/��Y�ƥ鯱�t�T�0>�.Z�W�������U/���b�3���`���@�[$����@e0!�O\��U-�Q�P��7���w���韺��t�t?��s\�D��zy.����a"�:��(J ������y��KK���׭��>ӡ
I	�mz���&���Q��ru��57��(�i��.��-�jVπ�T�M�j�þT�<j
�W��b¥6�E���?�$�WJ�Z��<r��N��a�m[���C�RhP&'�@�B�z���� �T�R��Y�F��|TY�$Z9٤�C�H�#�^�2 �U>��SBjW@Ou�f�8h�D���[PW8�3!־i7�T��Zk$��@|�)L��k.84�p=�[��S#m�}�*�5�����L�e�F�D�S3�i^p��R�-����'�)���ln;�ׅ`����2�c�J%�@�Fj�C�}�(�Y��l�;=R=|~?/lw��i'U��=]����J݂�3̼�[��)Q�X��0"	�k�P�b8!ghϮ���N-�H#
����������7R0D�T�bm˾���x��R|�@9�i�N9����;jw�y�����%�����-��BɃm��u.���`͠������P!$a��p$x�)#�cY�J 	��9�^]��ٌH���#��*�薹��.4�����"/�q-��<���p��&-���0�{ӁzkG�7NPz�t�q0��S0X�0��n��L�d��+����%V:���Dg �
m7Ȃ����
��m]>����x�aB�ܸ0U�=�ڞ�}yr�we(E,W`�2`/A�w�P�u�avC��Qc�5�bé4Ք�Ck]Z�b���L�����8VX� ���F����\�z��8�(�t�K,��{�)l��4)��;^Y�h�d�^���Y
*�L�2�4���̾;Bޯ��aŇ��i��"�dgf]���4"�}��[Q��Q�ͯ���s��ut�)��pGox��E�%mo�`��ۡ�c��D@���R ��
�Q�
\2��pb�M�z�ͪf�+��Պ1���r�ϖI{��[��N�>O�͔_.���5�<G�cb�V)���9BBZʽ��h�r�;1��
Y �,�����&�DW$�=n�������T���=%A��!���\+�}��++�tV�N6�����-
!��Y,�<���a�(ڹ�fb�����m��E�`����;y�̻��(�;e���}�~���T��=�&T�x�� ���Ɏ��|L�7wZ����|l�qR�<��S�]�Nx⊄�E��@�>}{��[w��M�����=B�ys�1���*Xue\�^܇j�(x~��v��(�&��PQkҐ����m!+7��ta��S��Qn�G���z�'���P��zQ���G�]f�Ժ��J_���$m��!iT��' ���8g�oH#g%/����l�)D0�$� d�f��zC�G��m!��:F��63�ҥ���'k�ި�_���-dkaP��e��R����ѧ��%�|ءK@��S'���m.N�K\���w�,���<b`t����z?[$\r���� �)�Ū��$���/�=��)��~7��L|P�
y�������6���:�����&�0��y(���[�v��O�0���J}�a�%�8d�g���|�׹���󍎽!��c�}�H+�	�/��]��ڸI�(8�ؖ�x��$2��}����)�?۵ �L��~�Y�kFH�d��V�VA�(��-� a\2����;�q�L�_��qp�x����V3�nىu)1]W�{��}���3�oH���k�튗ҁW�m��I�j��bq��{�R�D���}�.ǲ�����L��ۥ=�	���� ���in"w^LY�5$�F�B�\��6����\�S*��r���pG��s���+�i"Q�7{�ב����5��m�fh�'���Az�����ӏI5ݚ��̓1U���1�Tɇ�0�,�_�n��ZU�F��<	�y��KƊ�+�EC�L9���v7�}�MXJ��� � WG�)�ˑS�u�4��|-d�3�������b_A��xt!�ڲOݾ~��D��*��<1�l�`Y�s=������d.DuĚ΢� �ւsrȧ�4E��m�б��W�߈O#,W�cF#]lA��}���EMe;،DI�Koת@�_���`�D�	d���T�/�=8D��9�}l6bG|�`��H�����)��%B�g��٭Gs�/�� X% }/�2������)�54d���Zu[|`#"��ի�A�<�B�6��7�U~A:J��POK��k�{~ B�hug2/U>�������4�MPR�@Ji2(���%KkJ�
��C�sx8���_��KT/����'��!�S�`x{c�U�ՀI^���Z��4zZ��0.}�Wz�t<}���a���s���	�����,7���������[NN�G6�+&�l�{_cl������5����.������x���sh�^R�ӷ���j�nt�;m(��@�f��iRp�����"�����>ȓ����J �vm�w�ཛ�ʼ�7������  �[�V�s>7�')���Wj��]���nT�e9�5�3&�I����4��N���u&���}��GB`7���זּs?��U]�^�:��:��"��ݲ�fb�e1���rc4�kx��],:�4��AœS�ջ)����G�`6"B��6"��N��L�;�Z IQ�!�Iai�_�q
�kS+�Z�|i�g�f�G\�%�\�ۣϵ�h����m�&� �{p����~�'/�Cl�|v|��(ö{"{R}�O�8����x�B<a�
|-���bsD&:Y7t���,�E�������x0��x
�U9���LAM����5]@<��X����y��t��7�V�f6����c>��������X5�������#�|\��� Z�"�;KlD��Sa�z�*FTBjz�P� 7XЂ+�ĿCn-d��;fu/|�)�k��A��Y&i3$̦�A�Ԯsِ=N�A���w$�!�� ;yw�A�+8�o_n���Ã�ʝ̒�	�-�iL.*�LTjQ�U�	أ�7��j^@t{=��{N�n��T�,�l�U�Tj#N����^L`$(�Ê���W+�.�2��f��Vu�=c�|�}oD��˗7b�.li������3��z���M�E_*g�N���o-1������b� /h~9��I�ru��h���	�_־�
��f�a�U�d��+�SD��;����N@��ϝ��2�Ϣ���q>tm|Q�ʛWl����7�1�Bw�c�LM�I�v������ɇ����4�Cᴢ�Y�G_5�mD<I��!�*0v�$�|