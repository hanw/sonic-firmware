��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z�X�M�F^�@jaMz�����n��'�!��S�@�M��S��l�k�k+���R;}��:2��y�De��w5�/|{�{~��Pt���gOa�r����=.*��X�	u�Ԃp�n�hi��wB��{~�Irů�i���Ҿ�sc���,�ğ� �z���T����*�HV��u���iҳ ����#m�Q4w�k�)m�_��Q�����s���Ԁr��I�z��6a��|�g�#�p{�O��Fӻ���K�@�m��W������Ymg�UYp���_�}�"y�B661��0���<�-�7� �*tDI�C�;J��M�@�χ9�IRwz����~6HSE&�η�.D�T��o����MeB�ED� � b�?�k�,|����/������L�iXm`�Wy�5�R�z�Zp���$��U��_Ӈ3؀ꡉC$�u�����Ū�C�P8�啗��~$"7m��#8Zr����_G5�|�	k�"���?v������4>/_/Y2����wD �8َ�ᢽ�aե1���*!�1ȴ
��ۃ��J]�-��h,�J�����O�C�%��d�
n��F�3����|Q}1�z6y�������n��v�������է�e����y�9���|T�"}�t����'�Ų݋n� kr[�Fgm�l��՘�o�&!3��z�:ōQ,O�m�*鍶�A�̮�L2ϩ��j}�"⪒�A��ʬZ��BI��?lz�u'�7��Y�p���E##�,Ұ!�%���x�1W�>�`��$2�6h�<�3X1!��MDM�6m������Mh��p�[~�)�X�b_4:��Q�������I��#:�F�1l'B)�]\k�G:ME�e�ƀ��;�p���x��~QV�-��.#�E�*&ė�Ve�~2*��@����$�t�
V�W�CA x���W�_�S��m�Op}�����u��'Q�v��o��s��}Z�g.Q���YI�Vҳ�i#"> 4�c��v*9��X�f�UV��\HL�!A������;ke32d��O���~N��F0V$qV��p�Z��~�?7X!K��� ��9ʢf�!o�3�����bI����e��48��!���ѳ��C���D&���:t�� ����W���0=P�����۳W�m�	�ݞ���k2�{�R�j֔�T�S���hХ~�|<ƵzX^�xD}��@�W~,ğ^17���PDK�ȇ�/K�4���6�ty
}���H�����\���FӢ#1�ܤ) ��{�R�nh���9�m�^\��k�8�s&z�H#L�v������ZK�Gb��y�x1���_�y�Ӊ����_�q��ڢ1���k@�3�rF�u#H��HJ�zYO�	y���T��{�Kڃ��F3U���K^Zx�f�ppVO.|P�	e����2�*�O0����X��b18�8�xi��j��e��O�CI�I"3P��:�� �vZ��u��h�8�$���p}KVK�V?�����N�$g�%¸�{�P\�m����>k[u/o��|�op$'p&�����f��Г$���<$�m�r3A	=k͓�XY�����XI5T*#-M��BD�CC3-���4/��� ��K�J��&����$1Ak5
d�U�%X�	�o�-���X����?��.t_��	c�^� �UCY�8<�Cc����w����D�Ş$�ҷ���X�/�@6�oN�MA�3��Y5Mj�U�Z���m���9�F]��ؠ9��=dɫ���Ue���j׭U6�K��"���ţ�>�6:��0u�q����l�#�yp^���|86fn�����Ԃ7|n� A��*���JS��y�O��M��
���s�d����_d%����W�?p~κ{N?�(��X��1	����k��R�./��_��j�<�?@�e��z@!0�Jз^�2�܂�����;kk�6iăq�6<Xo;8��4�qA�L/W�n3��x^�����������m��]��"A��Ǖ���e����u
�Ƿ�,���ڍ�$c?%��:	c�3��P�gk�
��BdKIzT��t+�KY�0�:E>6(�(W�ɲ|�I��˲��a.q��p�bl�Bs�)��?IX���k+2Po�~7֙�`T=wW&L�� ��)d�èLRq��_L��O�_��܈����&C����$���ҿ�A�t���/���	��}K�Fz��k}D�N�xvA�i#��b�ۨHf0��0玊����k-�Sƿ_o`k�E�@0Hw{1Ku�W���Ȃ���Q����o�{Ud�/g�W0����z�U�u���g��JB�I�Q�S��O�Um瑾��c����&���	�v(H�bȳ2�zG��qs}�����l��t����C��Ҹc;�e�~��c7ȟK0VuN �3����]�W���O,��2˚'�Cr�^���C��K�W��v��=��,l�<������=^f�-����f_m �� �[�OjJ�7�kۀ���-`%�w�ߎ;�,5.�MG	.Q���\�=��իG\��f;���g�`�i���S���6�?+1�����B:�6�}�)�o��:�k��«���sĂwL�r�qA�[�^h�%��7vZ�7V������6�ԒS��
�h<[x>�=��;��~�g<#����br	��t��5�JX�H�J�O�K���E�B&�W�u@��	�InS�����`���A�'d+�����Xu�l����w��2�� ��ʋWy�8D���_���}�q	l�V	�il�U�t��Bf,�����!��N�����N��ϵu��)@��/�;Y�x,d�<m����Vf�o�9�����
��|ϫ�DH�G��'�,c���Re];�X��I�'p$�߇s���
o.�����G�jNHz(j�tţ��l�_Tp->��e�H�'��jhDyٯ�z����3>| ���P��Mvn6�V�p��Zv��ߣsAj��1/�������$���R>);i�b�.�GK��� L�J�36�N�U�����H��KO�{c.QDg_��P�ң��r���e�2`�r։�{/e����S^_����.Y�%�V2CEs �q�5v��1%!��-)9����ȋT~�/�tđb�{\,8�Dܥ�M iX��Ȗ�K:����3`�rB�Ҝ��+V�X�Z8lqa~b���T������x�	��b-�r�l�ӳ�n}'ŝ��B7�G����X���c��������9KI����LH�Us'#�o��c�����a@��=,{ţgR��.>�s�B���������n�KԤ�����iW�`.L�Ρ�-��\��}o��	�D�I�o:�����˺�K����{�/4*8�x��Of�Y@C��95����$�,|!E�%��������!Q>��셐 ��i���%=s[�,�=i�&���U:�nEc���$�&Ǐ��	�B`[	n����N�rB1��!�t1Af�~%���z2�Pj{rP��2U�-���<����dM��lҒ�X��׵w�V�KH�`�ރs�l7t��?�+Vb�=b�m��G��fτ��im�k'jz�����o����5#=��f:4ih������ʚ�� ��X�x�6�`	�� 8�&Q�]���5��06Z���7o?.Ih�er���7�W�˾'Fޅ��£�7��"dƲ�"S��x�����wɱ�ʏm�EfIR���p��5�(�d�ax$95Ň��[�~E�Y��¹ӳ��2e�W\���1�{�_�,�L���D��e7�c��.]�X��bjR���&���}IvL�7��*��<!�'55��^��&Kc,�M~J��*RF���t���4�9!�D>}F��w`�ޒ��R�����?�(ZG{�O��zO5��~Z���B̿��òc�.
  ����}&y�	rwA��k���V���=��Z{ο������5y���z��E��'}�gp@R��)�/����(;�����Zq�Ri��K�F�2�ۨ#��G���>;? ܔ�м�5|Z�m>�$^<�����!���s��/	�,�9�s+�l�r��!ThH-�#�O�w��5�o\EҞ���-�mFy���%lO�ZS�Z��R�����[	F��?�\O~8��x�1H����=R&%mm�r��;��8��k>����S��=��]O�&i��G!���>`��� �j]C��ꮄ.��FZ�N��������`��p���;���95%��#&]	����	�~i�8���4'�ǜ��d���q�H�M&�A��]�z����;6�B�Γ�̙b�J��,;E�/sW4�јF�Ta��/�w�!���i�V([�)R&!��b�b��#�w��t%���N튗m�Al�~+Z^�L^CFX�8c���^��J�*'�؂F5$(��;���;�zʁ���y��'�#Ř	i���Z���0�vܫ�	�}���qs�f�H��R0�}���	��/ן0VL� ��|.d����?ɕ%!Ji\I(0����]G7I���B�̩�_��d�>�BKkڒ�=+k�M6���}K��3������2P�줧=�5���a~«}���=��?����C隔��)�Ѡ����B&���jh�3*����t$c���4�WM��O���v�'H��Iʹ�>�;�b�0��)���DJM ��ap�)r�la�['P�m���ܑR�!ꈌc���/�T| A�T����	넆[y.K9Upl�)�7�� �N��J�i��R� �5�hl��iz��oLg�+߭�&��c�h�h�<?_�H�?���4SáC�*���~��]j�\��Q<�;b�����o�ߔ�܊��:��h�m�y|�O�n(Âp���\�?��~/�g�7T��u)��Sss��nv�|v�u��{&��MO	M�MR<�=�H�'+����$Q��8o��?&躧������zFT3���9v}w����9��0��) /W��V�<3R)����1	����Z���^߀I��qa�l��vJ�*$�~�	*qxfc��b�!���6�&w����ZY���L���a]}ܐeE�72'��g��%e���E�����Dܢ��(�3 ��2�rr��B��,�J�]bs�(i3n��CB���r�;�f�:V�:�k��L�"�����z=��MP+��[�#�ٸ����h�o�ٛ�9����s$��nߟ���Fw��F�L]n�dd �y�l@R����TkY��\��TE	�y^D�\[���&-�Ӟ�ǖ-:*:� bt����ߖ���[-RV/�@��̖�" /{ӳ��ƵԲX�݆{�����c$'�ϭ�0�m\��Bz{��2w	��iم������#�A�K�]L3\9�����*�'��2O��l��iX5��@�C�I,�����h��0��C�5(	z���M&vF��s�<�u�^5�CH������j��=���F{p�����5�� 
��N��o pp�ZW���g��G7��Gi̖3O��o63@��\#���C1U���rS����d�g��7������e�Qi�vA�n��
���C]�d��e����N��F��J�	�1������2��T��]:Ԣ{�h�[DG,���l�D����ܵx��g&$����v�6��T���ۊ�Km,#�e����	א�14�4] �#��>E��G���t�F8�����K��A<�H�U��ep揦���$�= )z$q7��{��d��Ҩ<\�@��|���̿���8�I��N>o�+�tu$
�e�U�U�*d�z%¨��
{53� �w�J��rV�]�"�� ?����<(��S[L��F�'��KY���ٮ��d��B��˜����~���A3��=Q�_L����W)v78��T���f����=6��Caτ/{���@�Q-L��wGo$���Z�/ޔ�u�8���$�t�<xÚtq����Ⱥ��Wn>�{l��Os��	X���M?�d4M��:8�M����S��8j�]v����1�kF���Q'�-�xS'����7���\9��.�G�����r��DA�+ղl��/�I�A�)�o���ӥ��f-8�Ѳ���ح�T�v�H����#��^�i�y����B{�-w3n���r���xĸ��d8.,~�U����-@���c͚z}|����j�-"�NE��HPs�y�	�
�<�6d�$$��g���Og^�؟���5�j�7h�?B�V���v�Y�r��ȇ��K����BVB��w>z"a/Ɗ�Rn������o�i���gD�_�V+�u � ��1��"�A�C_���x���N�\�-I,�$ϒ��6�.��;�v�&�\��Q�*%nNAПM��sZCՍ�����h��a�S.��A�i(�o�,Er���Y�Bk�Ce�����5xÃ*Y�<��i�X^
H�����HTs�X� �_�Q�݀F��w�1]��U����25:4-0ĶJ���Ӣ���7�k7���\_{$H<��Z�c�ٺeH��H�iۂ-h @̜�y�xg����8$<M=�����y�35��d���jq�0 R�儆D�k`��c�&<I�*�u7�3��q&�J�FO��~_u^����,ժ��	O��ش�������uDϽ(ɰ��dG���P��#��U��������-�S�^PV+�	`��
]I��\X��#��\����������m?�|m���H�	u�~�.T1.���?�q�%�;��!�T��.]�yL|���'u�T���l�VO1�ۻ�l�D���h�ӿ���7�kD�����:�J�f�Ϲvy���g�*NK}#G%�D#�}�L7��j�g��kh���D�ߊec���n:̹�9I�K��~
n�Z�4"���c�|:�n3�����P��đ�)X��;�P�W(SG�Q����~-�6��vk�	�]��ue����iqV�Z��(��5����9�U#���Gɜ���*�M�V�D�T�%��4]R(T��J��ֳ<�~�G8a�n�鴒�,�����n���|����Əo16@�}�ZS8�7�BGF��aД��~��ΧRy�ώe�@,=�"���:�KݱWK
PG��L�WȦ���c��������*�=y�^1���g+�=�[�Ǒn>*�K�O!`�笹�w�֛ �~�2�#e�	y?��GF��ȣY���$���N�RW���
��=Ȅ�bXO[�( 9���NA��pe�p��-=�XD�gԽ
._+� &i�C�ǎ��B���4=��k��O�U\+�$�W`���~B���Cj�l"ʿXO�6#Ćd>�f �":���Hc��ׂ礞$�qJ�8*K_���2`���.~R��J8��������S�M�V���G5��:P2J�A�r������A�G������-[���
FN�b�
��ޓ���KL�/Ͷ���V����\��z7�#W̑�i�;,z�����	Z����z��㺭._[f�����4p�+��|���>�%���m��|��	KEE^_�٭�t�� ���[Z��;L)�Ou�����X\���G8���c�z?���.*��ޭIK���I�ƺ�:`TZc� �GbKG�I�i>�����K���)����T�" �8�z^DTj,3����9k�V����y��uH�H�Jq��1⯌I�]X��ձ�Y:�@��m��贺�Dvn0ͣFH����bO7���D�?�Tˑ�ܒ�sAڰ�<�h���1�mήm�1vI��JF�Kp�q����m�K�g��>$��ov)Ug�Z�;Ψ{V� Ѻ�?�4Guyh
�{X?�D�f���ny���c�[�J��������3|����&:G69��݇^M��~�z�촩>{�p��L9e����4tq׭�S������-M*viN9�r�c8)]d�d�wn�޸N.Bd�}�9;"vѐ��3 Fm��h��O��ǽ��x>�Q�Ff��8M�i��B�*�����^��ݠbX���zT�跕�*�zU������y���=�|��e��6-<k@��7�O�l��-2�q�M������Jb��;�e�u���C$x�eu΂�6Ptgux%�9�1(o��w���h;�=Bc�'�j��aBv���Og����i�H#���am�Bg�l������֬�Gq��a�]�h�H^��T�J�Mv����E瑨k�t�i��33���,���9���*���PW�!ƿ:&@1ta0����J��1�JQ]|���Q5ҕa?9���>x��dr>�#�l*`b��C���c2�Am-if �{�s��u?dH�$=�㌍�x����ȌY!PF]�H��a�*�9�77�5z�cDل�KG�,cc�1��xI];���P">"O⹾4�xA�Dֻ�>�q��t&�_L/(�� ��d�g.wė-aq��ԳAO�.�z���'��S;f��S� X�q����v��������k��j��}��׿��)���E�����Lbz��aoY���ͱv��QQx�GFߜ�"w�sY��Z�����=� s?6��E%�5���u����E����'4���586>��!)���vp9�։���؀�e�C��M�/a9�+�-;��i,&�?�ߵz���¦_s��{3�[d]��ا�ƫ�`�A��=�LI�$��SŹ��l7�Rj��4/�
 ��P6汿�/Av��a8���_XT
@9j�*37����9�T8�ۍ�'��GZt��ƃ	қ=<9�wOԖ��i����g���u�uW�O{%��� �u
�y�,I��lp;}���٫����W!���n����ru�#3{^�jc�D�cR�*��S��D5�zV��\���5!���l�1:A��0���VoG|��?`7�R�H�	���5�bAb��;:l�Y|�	8*<�� �Z��@�����i^�ػQ�\{`����PQ�L�e� ���� �!�#RR��r/��vi�C�1��7z9kX�4y������v��*�V'�%�LI5������8L;��4��R^�qG���O.�6��<~��EOc���IJ��Q�Z�fXL6(��N�h1ˈ�H����՟��>����~ ��������4k'�Gq��L����JL��؋�c��6Zq3��i�*�)��;m8t3�r0Vhu�Ȓ�����n���p�� Da3e^�V��ЫU_��i����O�6k"e�wjlf@�w�$�%Kk��vF#f'��U�d��;���8�ts�E�f��2w���UL��;To<��_�a�tP���xq�X��
�եwZ*Dn�'=H��ی�J��t�2�y��5߁�$�/����o�]�{lk.�"�֡��0SB�g�,F�2�XTt9ZZ�H��#���`Ɔ)/�!��4-��_t̦��^F|(��#c�&�- ���f�m�NMzv�O�ei�t��*FgN�A/\�N����٪~�RE�
r.�k���{6�g6�vJ��4h2�/S(����ScL����@-�=����ch�r�r�����Ȝ���0�OO��TpU��\�NL`��n��l��XdSWB4$�u��qƇ����~Q�xO)f�Tt̒��CnPj�{���|I��Ȕ3N:K�ѢOC ��mIl��m�~$��z ҈�׻ww�҉�Ӯ��j�Y�lp�4W��skM��r�K焃�e�Y6D��3v��Զ�!���C)d?�����I@�*�[�/�ruKM�3�+~�*��&aJ�eb��d%iC)�ƴٱ:ćL�b����^���Z-����D�R��,8ǒ���m'���V���k�d�;�`S���37*�\��=�]�p�<`�;#A�b�\?=�L ������J(+{�qq�2$�(:�%}2�{̡�xɫ�ӧ=\MIXJЄk��H�Uv���4 _8���P����;�*�2d$Т��$a�*nH�������#}-@:}	ed�0*S�QR#�b�[-(H	O�D<N�J���A�zcqj��grB-��^��^䏲A=]GI�#�X�(��8+M��+*b���c�] 7��P����ni����Ѡ^?z�X{m��w�B4#f�^�u�]g���{��f8F{�#�c�bCЫ(��"'��G?4U���I�� <�������}o��l$�#ߺ�]�Y��R��VѦ������>�����XST��n��
	T,x^VUv�Z��);�h�S^	g��f�Uj3�Mb�a����ó��J�[����k%C)�ee���<����g��Z�N�xZ_Y�Pp�MR��N�����}/�oݍd�<��Kk�&���e"z{I�S���3Hʐ�=j�/��M���ȷ�c�ź5��ԝ�e�q]�֮�S�,��b`uS� v��
����A��&ϪEy�2��u�)��"*K����tS��� �6�]�x^i_����/sK51>�ٔA|�W��[Kmŉ�b�gD�c�ܒ�Uk�9�E[�䠳�C���C�eƒji\���c[���O[�q����c�K�es�")Fzѹw.�GHN�K��<��������m2*zTq`�B!�8������w�"ƇG���L,��Q8Ӻ �J�p��V���C\U�I�Y��bx��0G$N?�*^��:f��_K"�n{�Ӡ!�7RձD�Q����5 �Ԓ�+Sk�ٹS�42�2��a���U|'�4���h���$���~QG<oW���|e����[��*'�B7���+!2w�E��Tޒ!d�v+Ar	'<f�ݒ��y˝���U~��ϐ�������w�o��3g������? i8T֏�ы;k�v�v|?7Q�%�	���1j`B��!P����T�+�xu��?��^w�t�+�.�1���`_N�ޓ�p��n���������৵�����x[�Q�Xy�Fw�:}�Ѵ�4�aM�O��#��=��9O ͯ�Ibj�Y�YhI#��k�&|��]� ����p+ɩ��fA\������~=ٵ}�z8��r#Ծ4Xج��-�w5�J��Ng*t��x��C�0v�c�ﱊ���q�T���$�}[�I���`�lQxI޵vR�VM[r,����jxE�R����L[�6�I%(�Ý�7�M�ҧ-���h���7�)8-�@au��P��0� ������3J�8��
�iR�53B�x8c'�������[����WZ�>����<i��Nf ��҂�@�J�8E�6fR�`��@�c�4���r�Cu�O��~�5� D)����	қ �*�V��q���fW�O�*�A�^�$���0�[����$��F�{'�2�Q�E=T ���)���3���_��ϝF�b��0��?x+<����"Q�m!��&��U���=L�����	�X���4BȍsϮ"�B�o�[ª��}�\L���M�W.V�Oϧ�`�	I��@�>��D2L֬��a��x�ta��������-{��B��?�I�T��M��/PQ���D��`��U��'������:�{Wl�⦢D-�5-D��̡�p�h;V�����̇�(jܕ�˧�x �h#��c^7��$����
�����`Yzl���3�)�S���%@=Ƀ�����G���u/ͬ,~���s����O�2���2��}��֢êk5q���ޖ@���t�r�.��YZ�ЁR?�`;@y��-aM��ߟ�ExPr��޸�&���j�^E���Zs)(��hZ�â��u���3��VhLd)
���R~L
-�5��u%�Ku#"߬�Oi�&�*`	[h�v��ر�M9��a��üM��lq9�Q��6���97�ˈ++ �J��u�
��N��{�y�Rݷ�� T8�é�	�D|�\���f�-��܋�-ؓѡ����MY4{�~h2ae8�G5w*;=f��N�5ێ"dɎ9��:�x�����:Q��k�¾�g�R�5í������t�U�qK�M�/�<S��.�F�R����LC����=�	�pՠ{��Y3j�[�� �x�4;xn�d�P�2���cc:?��dG�G�sNӯ��z3�溳ܩ�?���y��=�������+�x׆��e9|S~Y(�s|�O�<m]zI���z�r>#H��ʩ�-���7�>�*����P��?	�"�RAQ'Xf��
�m��8l�́�^��t+���:�:L����2Z3��w���l$��9�Q�xӛ�(����i�����B�IS�g	K���g���k������aс��HF���`upԨR���w�?z�Vj��+J�pa��;���>��N:Շ��nn�R�3�q'�	'����Ȗ��;S6������!��{��5�X�KV�������.�0��,��x��z�~�1�`��kxO,D���"�w�;���Fa|^i�2�S�Lx�$�9=�+3����%���W\6_�A���	�[����1|�/��<����aߨ�Fy��������A=��!��J~$
+js�r"�2�v����t�<�"�ۧɡԽ�z;�!��l�ڍ�T�h�d�BM,N��{ǈ��Ē��_��рeHh��	�p�˰r�y
�\�D��"��'�����Ȗ<1;2�$R8VZ9��nS �vOC����Ƹӭ�|v!}�{���hb8���>�d=�K1��F-ӿ��!˂`.wM��<�IѤ@^	�C�7)_bX�\�]&�ޒ>_�i6�D�����n�V��t��0�-8��<�t�s�_�Rt��m�y){���NO�U�� ��ƥ0c|�qᏄ10Ta[� ȡἊ\�%ц{�f8��(�䍂(��>����v�1�n"6��Ņ�_�3�����7��7���������b5�OÏ�d�O ~�T� =��6dRz,��b�q�q��m%?��\������H������s o,e���LZ�I*W(�/������#�W�&�6E�|C�`��9|��M��B��)�)�*zx��P�B��u�LA���Ϡ���}�L1��M�s�~*��ѳZB�pͰ�Ǟ��x�/�Ϯ��V�kN~��=�����f��t�=&�����ہQ�:*������wO�v\a��\N���HS�d���kn<�	"��4 b�qQH<8��1.	ID���c��}r>�8���AVV/C�1ĭޚ��u�1:5z��XH�4��aR�X�>1Wy5j]&�6�ZI^��ӂ8bց~�u/�\W�X�A �c�����~�A��'��=uN���u�g�D��"���|Ҭg'&�J%'s����g�(+;)��,������'����	h|/:a��7��Z8�A�����}�\톪�3��(,��E@�˙m��Aң �����{��L�Ml���69��[��R��2h��p�7�z�qKu��7�4��/H���2�'(��k�>-��k�"������!��6�K�2U�/����LS�,׺�N�������y��ܿU��߂��^KG�?1��~ �V�'�i*��f���� ����xT�>�)l�_��&�����K��I�kڇ�������g�CZ+48�$�y����xr��-����V�0����*�������͊b ��!� �_;ꀶ� SU�GU/S^d��A�/'�D��;�,��54��{w���u�P�&;�H��uupR��KM7��+m 4�e0�y�dq��8��D!�ù�[Ԁ�u/�X�Lh����V����0|q5iT��X*?���9[xb�`��Ĉ��2&8�g�Ǩ��mD'e��U�|���,gT�	�\�il�?@�0��Zl�A/�U������Q���:P�+!�V5BJ����f�;��44����K>���mA���oeu5��:��:Qs ��@��j%�\3Oh���s��#��䛮��-5������ȡ��D���Ú���jP��6��.Zg�M:aYc�cL��g��77��p�睞|����󵬾�?��/� �u�)�V����DBZи�!����2�m�Cǚ����%�t�w�2�[[���26xV��s�/��
���y�ˑs_����S���;�}%��AGc3�R!��g���x؂[�I�S'�,��)J�&��c��I��ձNM�KElpT"g(v�u�Gؠ���֦���� |yͽ���l�w&��E��)�\�s`.��Y+A��h�l"��5�Z�y(S@\B��2rכ�gGț ��-c�A������3���N;3HaQ��˓�6S�����c��3���r,rj$҆D�_K�c�z7�G�5xU��Im������k	���'�/��"� �=��ՍA�nG1�a*���7m��A�3/�W���a/NK��:GѦ		f����݋F�͠�w�����������,q��e@#$˯78����Ϫk������KZ�m@P�&�x�y��:���
P:� �o�(exe9��lК[h�@�^���U��X�iFIyS�k�Y?"Fַ��u� �ֹ����}�u�����9:�\}���M�V��(( �3���V��4�Rx
��x�R`���ǥ�BТ���Q�kQY!y( #�F�?�W	�����HE��o��!5(��!�q�?^����1��D,%�N�ь���N ��A�խ����Ћc(-5���]�J!`�vA�[w�xj���fz[��"�7�ޮ���6.�������G&�<x���Y��՞�j93kk��(��w�Vjq��i[�s�3TJmM0VM��l�Q���9F�}���wk�\�=o�u�韔�2�,�:X���+$šI��`p]P�$z��-x�)&�3%��[:@.Ο����xz�+f��.���Y��S��F9K���"�l��	5��A�� 䍋�:�WP���2ʲ�5r�h^fݘ�A���G�~"��5hUVY�h����
�M��px�gwD�"-7�hț�+�r�K'Ǜ5�)�&x&��T�d����v� �$<���!�'��)�|�SZX8b+Ç(]eж�X� ��t��2|�9(ě�ʶNO�8[Ig/%u�#	��`1���H��0�)�����9KΫ�0T4�EK�~M_a�B0In48��{?�[�'��¬����{�E�O'{�������y�u�bQR���mw����1�}����T��YT=��s�`V,�ULg���P�q|X#R`ӯ(�[=45�P��]	j�9p�s�.��ι)�J��1�+s�mpuv���qw�g��>�Y�(��~�|�C)��hq��Z�<G8�G�;5���D5C������)�r�Ua��@G��K\�ȠdN1� ��
&]N)�4�LR���\���y(�G���Ќ��}}�Յbw�̤ Ff�4�X�L4Z�</P��]���k����(�o&�e�W���	������i�6�8H(����%?��[���XΡ�����Yv�x�U����bP�!�Tc��Hl`�$�%�e�tp2����2yh�wst�E6|��dy\�0�t�D���n	&T��Ex���r��F:������ږE�2�`��z��>OMf��\	6�4��M�r�ć�vpIn]��ܳ��Nf��ĺ����3lo2�-���@�=.��<�s�� �M�
�Hе�S�W����Py�d�F��0�R��*/_�[y
j�&جp�f���|/1�?�h�N$b�)�rF�����TYC�����	ɪRR��ȟ�̊�n�rp�)I|�2ˇ��Ӳ�ք���(4�(Ƣ��{a��s�ڇ�	�2���-y��u�`�I͋��		��~0͒;��w;9���3r���#��d+��زp�V�6#N��~��1��_�H�2�7@ Q�<������ʪ�&���%�;m�~4�|!��p��Z����igdY4���[OL�)�8+�v�{�A�T˪#d�h��.ߢ�~�d������H��f/dډ}!��Њ��@�)��<���>T��N�} ���r�;�i �Ѵ�Zԥ�C�Ѓ�~�׾K"�G>��;)����cb�V�F��uS�	�+T�>ο�������闪�,��ݢS	1dAy���pH4sbxX)�u<D��䀢��"�:\'�*i���ܱ�Z,O���+�V\Q/��H��v#}��}�����D�m&F�l?�����f��I!(N�H�@J��͛A�9d'�?�W��ZO�}P��6,KG�:�Z���LĂ3���a�	��C��hG �p���etƺ&�����(���k�rޭC+�Kh֩:���/튏\�̭ΊȚcp�	Qqz�H�
�4PրX�Ц�@���By�sa)W7�4��w����Mcp�	>c����1S�}j�P$�Cs���:�|��:����������l.��.(j��O�*���L˓D���ח 9���{S�4�*
"�+����(���k �)y0s1e�i��<!~?�YC��b��u��O�Xm�$#�9�}[{�J_�!%�R���oT��>��WwW`'C�g���������Yb�j�B]%鳽7R�+�v;�K�A�+ٲ=�@�CyE��V0�U���4N�_�T#!r���A) ����Hun�o�0*��e}�[�Z����Z%��F�WE�q��Jw
���g��B�1S�~,K�����о�G9��&�hr�y�����������{c��˓7ar�vb��Җ��.��j"q�ӌ�r�����ι�|S��z4����ǥ伢2����ƹ0�pG���^R�K�ì���|w�c�;�VI�:V_��S�Bk^;B�W������
��� ��w�%�f���L`����I3�Qό(���N��zw\���E0����)x�#�%��GI:��9�Ґ8^0Qg"����c�!���.ah���1�2:�����V/o+��`t�y��X����TДT������nȍ6��eҧ�L��Q;����Eڑ�<kq�]��#�3%d)cW���m2�LR��53������4p�q��c���1E�"�	A}���d+f$�g����O���w�n}�X�	���0�YdD:S���=��ΰ3N�����x�,�Eܯ۩�Q����7��>G���y�F	�%o��xJɑ����WK���J�/�=Z�b�rKA��\�Og:�.Z�O�h�6:������1�v�7���txS`[��#D�p�wLjV��
���;��g6W?��C�75	�0!~wc_m!_������>�-��͒��| ��1 32ȹ*y!��N+8����Ԅ
;��L)wd�OFH�I,`�_p;����Y�;1�z,"%[�.�� r���o�O��5B2:��1��"�\C3��l,���I�(1sf��_��2�IM�[n��`���ї~&��̉���2=n�L��K�0w��Y��<��
a������C���G�B��g�)��ꋥ�lp�P����ݹ����;��F#���]�C
+c4�IB`�'O�Џ���("Fp�*��zKڹ&�Orm@0M8�C�lW����[ŧL����,!����{e=�,O����I��X�>3��H�>~��r}����}Ӽ9Xg�֘k�*i��#��3��O�}�Ci���M�g=�ڸ�^5<��ђ�؞Y�ŭ�
)P$����������_��_CżOm
>C��#o��s��������>D䛥��*v_��r��9�G��]dO"
����%uKDNe%tť�/��)�4�����;tc'v2��W�mQ��{#�
΁��S����Knb6XG��$�F��n�2�����<�qmB�MÕ�xY�w��3���|��x8q�?u@p�S�2z�����2)_���r_�D}e����l�GY��=M5��y�7>)�K������og��jz��]�q0�ߺ�D��&*䩶πN�z�W}
�0���4.�j��>i,!m�,࢓�V���B<�A�3R�Ea��������^-��l$�B����si��f�w�g9Q��>$=,�奾#Va����W�;9�1���x8}��X��n���șZ�_�;Dl��S)�?�د{d�e� |Ȟ��b}���I@&.��W_Y*���/�k����\���IS�x�X�hf�euQ�Ö�p��Q�yE�r��@�wx�H,(>�{\�\\�b؍G)5�l�����s�h?��[�	����%��"����E�$�b�>,�����ع� �d�%(S���������c����n�B{pTP�~��X��� �6�2R�����"	��O�9{27�Ŵk"��ߑ�,�k�@��9��������^�XȂL ��1�e��C�l�<�	S%�=����<��%����;Π.K&h�`<�eV\�(e�':N?��p�ZOu#�S٥�T�R�*7B��R��C7���r����C�±`TC7�f)3U��V����=_�cL�E3`�������<Kp�X��"����&x��\��_`"cB�+DW�付Z������`,�صw�'�&gf�eBj����k�a2�]x���')c��D�kI���.�SDvE�AHw�
�jA���(-/��sT�#L��]h������L�m"���ǼNۏ+3��>L/���;����|���R�D�V�xY0��A��v�Nٔs��W( �/?%���*�V�e�w��L�m���C#Fl��d������\-��K�\%	J�Y`(������=㱺FS��i~7��x�v�*�|�H�5����T�_ �p<{�u�?�Ϻt]�D�o��0mf:ul�=u��Y�mi�R�XmsMG�K��CWPzQH�J�Wot�~���, )�@�`��Hy^���f��^�A7	&�*T���N�9L�}M�k*/�-����+��GXu��Q�n?=X�Q9��j  t�����S3n:�^����Br�)�NSR��+��v�������#��b/�a'
�F��>��T�a�"/�o��	�h�g�y�*2�K�	�~]��hm^�X��B�����R(���J,�mU�(��i<;Co�"��ЭV!Y���c~p�E&�h�˜\����(S�@b#�v�k=\f�_8��4�����Wii�2/��q&
��������4&�LDp`��
�TS��$�e<l����[p�p��Y���b̗��P=?(ɓm��틑�@s�T�l��ǏPf�Ւ&8��S�e_
�Knʹ��(�,��"?�"��ɘ��ͅ�W�2!K鵷0NYjs��7tϨ�ц8�Tq��mGg���[m�ه�>י��,��t��bfR�\9�12qL�L�"�1˭䯕�.�+�O�	�� 
lG��	t���q""�E2��.�5L�X�r�V��.Y�p)%sR:�8��H׻��V�)�������YM�:�����C��V�y$�����k0�GP*��H7�3�?
���b���TdP���z��j�oB"3��u�,m^�H����X��?�w�s/�e��|�;�@�FI�ܳ%�/V��`Ϩ2�����mպ�����)�E�X�̩f.��Aj�SHNLR��jW�M���.{g�/��i���8G�K��˭2�h�z.��e��O���)q2���6�/ci�7��#S6)�Z���K��~�a�X4�ꤵ�P�ϙUHE� ��R�'��u����'f�u^��\�=d�ں{�%F x��o�|E���.k(م�Q�$�Nf^ç�UN1���~魛TK�7� |�[Dt�c���f4�b-,gA4���zp�f���e�0�I���{C�֝l:�k��ܟnU�g�w������|_� �ntS�5�?J'��
���R<n�
@�T_q�y���E������=���V�����¢Y�����^,Űxw�,j�
;܈�ç�7�kZ�˞�/ϊPَw�B{��q�L4�V�	:+ۻ&��@OF�|Lt�o�r�=�|�X����F1�1ݕ�?-R���;����R)[�Ѵ�s1"o�3�HWF��ڲ�ѿ���<^�C�t�A�.�O[���|��3/����Ǭl��W�j�p2�n=��V��Pe���f�����	��������q#^?�\5{z��6���d(���M�榒̴�V��qÇ�{h8BWa9b~�x��c��J+�<�s���"�C�>%��"p�菕�]���8ǻ/���&���׬������,¯EA�f&�TJm�k�<�Qw��<�=CB�Q*��;�����/��j�v�N���z�{ϧ�ŀ?㾓�u��q"�׈�A�(�=E��E�.�;����ً>�s��rZdON�8Uw��h�{�\�rǠ�q����Q��Sn;�w����z'��T�%"��(�GP_�ə�8[3�����:;?R�C���R:���p����_Z�4gt��|_g1G��H-�K	#�]��>�?x��\��"�Ga��N�
>��� �I��MsU����1����1���f��P~��Rc$�����_�W��/� 1�Ie�	�J��*�"�jYUV�gs>X���Mg��ԣ$����)̧�H
�!U�[��}W)��򀨿��\B>���zdٲ�G<��͊����K6;����	������v��)����/x��k�˻�3�u%������!�/��X�I8Fyu��� �6���|������#W��u,�����X ��(8r�#���)������#��X.�*��S�!�NM(,�w�$��ǂ��@���e �v}7P6n��ՠ�"���`lLb��ϻu�o��p��x�önY��q�6�.������v���C�͇�ے�}���r����������`'�>�s>-����{s
���{`+H%f�� T{`�M{F.��A�TyX���̈́��gU�@ fd����V�dD�|��e�=��j��K��][����� ���`����)��=���h��A���n�.s�TP�4R@P,)(��daN&,�L&�O��;�|Q��[n�ʞx%DѢ��B�ڦ��f�({���:C�������h���t���Սj0�?���#�ahpQ#��k�c#����A����ȩp�����)�>�D^U8�k	ܷ�������*J�dA��t��_D��k���� q_���L>��r�^糈ث,>uW�~��{���5��YX��9ͬ ��C_��煦V5N���T�����KD-!Z��&����-�j^U"�?�ѣ�{���Y
���E�єխR�ӣ������̎��4�aV�>���~���u	�}�Ht"���0՛�F������ ;�������g��,jҀ��*������@F"�J!�}Pd|��9�[�1��I�����W���\ZG��g{�������}0a�I47�.���M�z�����Y�%_}�o ǅ��@e7?j:ݺ"�w,|V��!Z��U'����%�i(�g7h3\��n����	�։(�R��$z@���Z���/�;�?��[�%��s	�����_�$��R^��9M/�}J>���|��o�`95!nCCX�m&dm�G���:��NT��b�$_۟d�Fp��m$�c,Ï�K�Ph�-���`5���po	�*	�OLHuL؏H�=I�|)���E{�ɀ/�����fs��NW�!ĉ%<�^XOц[z+k���B�wnJ6�
��cM��#Ynjw�����2�d5�B��"Jh��%-�P�3Y���a7�gDS���h�������Ô��-2{LKF3�k�9��'���w���S������?�+�7�>1�~V�-;Pd�����i��.Z�jWq܌h�(�ͻ~[���@�m&�^��2�ΐrr��R$���b�͸�%���4�|r&fȬ��99C _x��&����'\f��y�.ww�5`\��!�����e�I�G�j����3Q$>�g�Bh��E��	7%vr'�Ӕ<ˋvI@i�c�NS�j��\z������QpnrZv�Ě�'<A\#��jVo��}��?���?���Q�HT���B$!x���n�)���lA�nbS'���ӊIF&���<E[{�f� )��~�����ҍ�D�{K�k��w�K�rJ
B�8e�����o���n�j�v)������'�[�p�H�ϱ��I��������ҝ����d�ͷSs�T4:z��牶��3GL����1Zd��延W�6��
Or�>#2�)�c*ԿNֹ0"�GX����/7�Խ�v�[߿̈�w�a�?���xˬpUX� u��mT2��M�"�W^M'ེu�>��Wנ7cֆ���`y��?�X���0�C��:�z�(x�l��y	 �Ta��D`��I3+�b�^Fk5�C� *�RF84�3<X�>l�/��|�q>�5�J̨�uT���Q������j2���>@���a,��`��q�i��-��,W[�	lϲ��&?��{�����X�>S<@c���n~�?ϼv]�5��J�B!��p�ד��f�ft�*&o���6+7�h��%ELΩ�T�@:3+1J�*��7��N��W.����C�ޒ�a����.S7n��b����:�?��2�p�V����+�vj���T.?
�%�} �%�$�ڏΌ'_�^O��|^ �o�"�d=�N�H+ZΚ�i�k�������Hs���YP-�^������ܫ��P��ފ��X���cv�%����J�t�����~T���t)x��h7q�h��7�~/�����qi�p�Aj�:`ڱ��a�J�Ka5L4/�`ug�gL��|$�� ��΃���B > ޝ����3
��Y߃��������/�0�YY� Ӓ�wRnG�hHR_�i*+Ǻb/�@҃�'��N.����(j�l)�U�Y'�4e�C���k�K�/�Zp�gÉTB�{��Ga\�N��1RӚr�HI1�3��}FM��)o�M���7*~�oYV0�kg���	��d���&J�9�2�ϒ΄���ذ���LV)>�U%�	����;Q��,�np��,��Ỷv��o,P�YGT�뽖��0��0Y������%�*E��"ŏ�����w���Sw#�!�hRN���P:�X$���'��b� O�\m��k�sٙ3	�c�\,���3~^A���bH��5�	h*q����y#1��4�l�	\t���}7��Q��2���0{��K,䨞IF�H8}�֛���1�4I;"��M�8-
���]�4��d��~T"C���I���V��<�_��2�Fj���]�1��DX�T��fD3	�-�I,�ق�-�
Ż�^:,7�C��|��������c��$�D
Z���A[ɐR^5�ֳ���i�ӡ*B��^U� Җ�K��y�s*g�T���;��e���^�_�O���?� �M��Ģ�+%�� I�x���^� ��GD�Bm1Nj���K����C'�:�