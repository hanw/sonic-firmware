��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z��K���v���U��3̳f+�n�,����'о�P:�����u$?�b�Em>TѢ�C�I&�(�\qlw���|��l@�L ޶�2�i*!�k��S�y�U5=Ĳ����'��N��킃���#c�TIq�o�ICJ�r�'F2�e�B��{�o����u��4�.�36(�h��a���h��цj�v�{q�wN��J���ӽ9q�g�������WI��}�8l��+�曇
 �v�F�I`"�9&�(�.�-�m������P3��Z	����|
EE� ���:�;�H��n��Ohmu-�d������9�޿��O�a���t����!p���T1�ν���Sx{�`b�2E��	�	������3#k�y��P����i��-,y��L^X�W�����������݁�goto[���-����0y�-Z9Aɬ�v��iGq��o���^�l�z{���b�T��wߧ�P��֍��j��%ڕ02�2�|������dI'��PHV\����=t�5� qX�����ai'��6O�H�����(��fo-��s���RH2FI��?ʨ��p��:�;kE�9�+���Qv��Q��'��U����w������E�\�������)�B�L���w�>�����aH:�|F��
�b�� c<_�߹��e�^�KQᦤ�cy��1t���ȱ_�c�Vd�����ji��R,& ��*�����J��/�i�8��cT]p4�L����6�au��DAnȍ��gK�Պ��	���	F�5Ȣ���%j�^J�;?�3���'�������.�_�]Y��_�t�9�Q�'`þW��i�[	�W9�b�	�A4�o����sk���� ��y�
��*��D��-����p��L��ؕ~�o,Ɏ����O�owj�rg�6<g�V�{���&P56Fl;�_�G���V
���C�_Qp1hE9kr(ӯ�_@!x���l���2Q/�K"@k?ڮ����p�@����,u�+R�����,�*�:���a�h��0~@�~���8?��G�T�
�s�Ht��m������zS��E'�sM��v����)6�t4T�?��.�{�*��xy6VPe#����5��A�W��m��;���؀Ѭ��yZs|����Q�A�%E�>��A:��O#Q��N�{w.ʤDa�ېE���\�p����^BZ�����y�E�
�E6�MA>���r�^��ED��2��w�kR�{<_��-P�#}�� �[����B1�߹��H����󙋲|�%�[F��?q:�q��9�H�D�yF�b�U�&�&9H�y�����Ck��l��:��4����H7��ߋH�((�vr�j��Jڌ��u]����m}p�
�E�8��CAƱ�k��} ��ScN��ҽ�4b;[!$�R���˟~��Z�ђ'/j��&
�m���M��&ƃ�Dl[��f��a��5�ߵPPzE���d[�;[���+U�����SR�� ����Z�@s�C�Y���8�����X�G&�n��.�lW����I'R3x'�J� ���q�[��K��l����O��e�]V=4A�\%.�o����I:���՜�jBwi�������_ĺDoc�$�7�ʠ�D��E������5���X��+Zp�ϝ9���'�M�S�W���kS��F]��oՈ��i�>G^����s�	� [�T�$�d<�e�	���:c�5v�(���x�̤=+i������"�Lĸk9���a�J�у�6��1�� �2�ېC �4���/ԒM����wFL�.��C�u�B2�3��/;:�̛*�B��˲�缪�5)VL˚�[-�R���	D3n�X�{�&��*��G	tB��M5C&�j�dEx&O��E�����л����؀��d��9�rKtxT�];�N����[�]����t�4Q�9�x��@
)�ZQ�|0h�c[]i�h������)1|޳=Y~�e"� }^HB�j}m�@[0�0�4�v1,L�f�q��}!8٦��C3AD2��TTƤ�׳1�[W���y��m��Z@�6'�(Tp�_ξf��O�KJ���E��(��Y��Yd웁R�R	����_�b0���D��}��}Yj��`�{^�q�\$���~���4�-����A�H����`�-�}�KP��sX�":���!ꮚ<޺c!�j�� u�/L��������I�C��!P�����a�����L֥���
7x7�����F�E����̟����ڋ�@�����/�}뮟�E]j5�gqϪ��̃�;�P��J�����g�s�6ܭ��[w�/�^�t\*�1ƣj}ѕ�kT;�A�#���_$��s}��y�V�
;*:�8�U���$�ړ��VQ�����]�s�˞��ɹ-�j���@��퐰��6���\��o����XX+v����w$�Oo>�)���Fx������(��}F���rܡ"lO Wݣ�Fm�ji��e~���}&�iK3�-����������\`���
��Wq�@�a64^<��P���H�<���୆��?���O�N��c�����W��S�J3����,�I���^�҂jH�n���.��N�{
���h�P�S���g�~�E@�׈�~��
u$D!����fi�R׷]'~VA1����Gی��ꈲi�f�e��u(Z��zi��������B�ף�/D�z(&��>(3��X��Sآ��Xe�Y����,�u?Lp�?�����Y�N�f;�I�tmo�%2��r�]��y�)����`��	� .��
A�����s�������YC-'?\53��/RZ���ʢ���`�v�i:0)����2����lL����%�����$R����@'=�3Ⱦ�$_�ĩ��g��mZ�I�Stt�@�D���^��HOX���)����.��v�)	���!t�/݅�b@rr�w>����/�3�㦊������P�����[3\��t�Q"1�E'�U�����V���H@�#0ɩ����Lj'n�TK�D3�X0�t�N�o��nO��0���C�u���r����%A���h�S�mC0GP�ys����i�}�Mv$����#9\��#
��� ����?�K�z�Q#p�Q��	!�(ct��T�=�A�Y����0�9�&��ZC
��P�N9�\øد�u���8D;��
r��q����O�%6��S��!��H�b��;ñ .�/��OI>n�k� ���d�S���fR��oH���˹�����\V�@OR�r��|��+��0�Z`Q
��?`-�yc��H�#�l%8m�qe���4{S,���y�X�@��.W?�j>n���g��0W9c�� ˺;1QH���8Oo�ʑ�����%SS���'Ag���Ä��M��k���enK�@;�	����dJ/_U3�C��aU[��'��D:j1:9�^�a49������pN�l�A D�^���=�3������K����O,����-�t��=��C����AL�``�G��ߜGey�1d,UI�mq}�))�Kx����j����F�E���
���� }u�t&�e�w�,,�1��>O�0c��CqE�����@��އ�*+8J��2��R�%Xq��Z�|ϳ_�ej�~�L�I� ynM�-�E���Z$[(�Y�z�����I;��-����}�\�������A����4r��	���%v8mu�Dd�J��ʔʋR�G�RtfZ�9��-�v}���PE��\�s���=������EU$�?V�)(�9Ӎ��[���[-�Nx���l�S4�!M1�[bJ�X�I�4��v�*c9൵nPP�j��nыvսN"&-�4��K"�u
�;OWY�H����>����#�{�g�7M�&,S:��	���$O�rx�
k0���cF1��Y�>eu+?-l�ډ�J"=K���i�iza��%sYH5��XAv(0��P��H�@~g��T�hQ�V��ʌUs����p��מ������#^ҳ�Q
AKtF:�
uB�����	�����EH����)����'���?�Q���A] ���T����'-в�G`�qE	  ���yY�_j�a�:���
�pD��E9�@OQS0l��nN�މ�K��IE�ڻ�W��T�5�.PCo��Z��'��t������
g�,fB��X�b �P���5���>�" }3��D�q4�ٺ(	���p�����z�&W�sy�2]<��T���>D��Ul����u M�	+IE/o�އn ��s�0�0��ٴC@&T��� U�LUOћ�l�ں���8�!.�=�u��s)%�~�m����y�	b˥�/��4�Xos��[K�F��]�Q��
�\�6fN",Y��bt��@�3t4�ԓK���_?�yS��g��mkE�h���,�/
l�9=2`
ѯ\�{���C�;;ң��.#<&���a��"Q��	4�[��_6�9��0	��C��qӓt٪��a��
�`ؙZRMlZ�p1�:���$�����Ӂz�CG������'R�N��t|���a�vߡ�����������H��BO����pn�|��$ �i=�}��\��e�u��Vu����+��;0+?�Ǔ��/�Qe���"�rMx3#Ϲfح�6+�~�'������7O�j���	�B}Y�!Ut���҆�V�``+�a޴
[� 7��	a�<�;�F�r^XMQ�ª�/�KMB�K�7�"�c��D��ԛ����ys F����06M�yw�?:ww�xU͋u99,^�L��c�`�#�7�� �Xާ~O��
S���&�"����;^C�x1��uӨ�2�(�ߢ�|	2h^:�����|7P72ĵ�����*�K]4"�v�(n�q��<5���|`帍�s��C��^V���aPx����;�T�V���ʨ���.3�{�-Y�#٥8`�y���$ �U�ZHCߠ��T_�2��R4��/^��~��B�?�i�L_A��łY����D��5>��]�w:��D��<���K�db�|�*��=�Jf��?�S�Yʯ�Z&phIA�Q{ T��/t�̲��	A���0����8H�.�8:��7v .6z?�@�p��3��aa��@)@&���a!��6��C&��)�\0G	[�% �#�Z�{| tx�G��[�j�<G�iu�-��5�X�ky��֧�(�s����&�����@���������,�!������%��".u��N0�0�-{����
Jh��7�+~���w��7�&���mռm�Z�Jx�H�Hz�Ha�4�Ͱ}��H�£����1��:n��#ջ���P�����m�%<�՝4pE�>�ҝ,��*����j������rD�-˰��nw9,�>�O��XlF�� �dv`Z�[�L����S{��<T�'�%�2������������M�����\{�T�/�9�n�$�9U e>��zت|������	��t���������IjS���oua"'��dmU	A�[L"��V�v������(���������!������E�Ț(�$Β�G"$�克��R�6h�*B�tٽ]�nL=�g�x���v�KMR_wƂQ�*´cP���Q]V����������QC�m���>�7-���R+���_���6<��l�薁��G��!g�nO���G9R��Vw`�px�(��)eO��1�xa��$ {�F҉�h2��ӝԭ���l�nŐk��F1ܠ؇zT��aWӹ��]�(Z�k-~b��rr��"8*�2���	����*�i��cЛ��>���P�IB�(�21�6��T��q��z2�(]D�@�DM�	�G���Q�o}��M^"���o(�+�k�~1�;�X֗�i.������HDQ�$M�G��̈Or�2.��=0�>YP])n��c����NN��n�硢)}3Bd�h6D��-�`���M���v��N�k�[���$��r��\��I�AF��-"1���B���A���o���hbՅ��*���R"mU����j�C�!S�[7�T���EmpO���IZ�qW���@^��v��B��+Gf��.����9�����i^M��EMjA����HP��U"����$�
si�!'��v���&�;!!,��]~�W�����a�S�_x�)_�M�9�\�C�X�BX;�F���Br+�~L�������S.� ���!��T���'���ۃ!WJ�^OL�B?��N�F(2Yۦ�sff��߅@�ć��N�Vޝi4[��)�Y7Oef;pAv�/�	%�|�j��WV���v��6����t�PZ�6.���!��Ҍ�hU��)��6���*�M��ʞ�B��f��ND7�)[�o�H	W�A�[J��f��ȭ���bAC�[L2�(u����z�/{A��{K�=!��G�������<�ͩ��%�~&�7H?{�1�ڋ�������(���J-XO	:�
o(��VL4�A�8u�6���î:ݷ=sbße���'�:�y~T���=2�^z佸�اC����[ܙ�ѾMR��>U�v-K��W�禝S=�>�q��޳��ر�_�ȤK�~Pb�W�ᴯk�U5��pƥ��������o�aKޟ�{�V�/%�%�8�d���i�X�W��dU��Fџ��ЛC����R�qn��xv	zr4�ʤsK��;�R��9��2h<���^��� <WW��Д��8�^���5��X��_��HZ�3��š�1�"?ꨴa5p&�m��
��Z�Ok�1��+��&�}aZ�		<s!�ɼ���k����0����e�\;��B��%��qi}'UR��qZ,,@��ڕOO�A��}P�Rt�����^Z1@M����j���;o��VH���"�7�b�=J���.��!���Kb6�~N���%r����(l�C�u�0��tĊ�܃����r����}JU�u%�9b�~�ޕ>5��QZg�5�\lx �X�Nv>�A��ᱨ��Q�t��O��z^��TE^r ū�J4�Fp���$C�	H̸�(B}�I��5I5���uj�E�^�j,ٴ�V -�n�s�T�b�(�I�`Y���N�n�׉�6y�|��]It6�p�z q{��y�З
����'�5y$�*�v�P�i�I�T��m
���VGd�	ҟ����Uخ	1�41tY~�5�6�`c<yH��N�FEF���Lİ[t��'���I�3M%�����*=�`��n�����	���5S�9~Q��ga8�y��3�]N��@XO+ Dg�{�$�����鋏ؐ�X�K�����o��ܴv��������s�5Ϭ�����p9Z�+"kv���1��S�ˢ��:��:�j\s�'�`�骦4���̽N�E^C�Cݚ_g_u�~�U-��f.��Nm���d��>�N��'���e�8�R��S�̂Q��Z�x��wQ��<<������f	B>�!?�`-``l�bP�*�{m@����_DU���`��v�E5#{x(.azV�*�����*-��ԭ�;�[3�ٛwC��㛊wf��T8���P�]����0�F$�[�¾���@F�IVz2�OW!�9<	�	b��)���҆<3�>;� mW,�<������'w8��Wctz�)��6)2�+�Li�Eu�-T���6�eI���C��o��h!T3;a��:�y�oQ��fdk�t���OAlx�2K#���eb��D�#���&>.�6W��<>��^i��'�������z��{A{���ch��A`<�7P�KT�z"�ܤ�뾥�0	��eg�ltհ���C�.��\V�(�� ط.U��l|;_�����7�m��1�4N�Lh�~-�a�X\G��n�P �����(�x�g+��g[ �BWÑj�텸�� aȱ���C�N.�y����Y�5}m�;"�l^u�g�J|H��D�U�OJqDd.�m�ou��?mաi�♂�����d�=��j?�������2�RK��Y�Cd����q7Wc��a¿�ў�c�j��݀�ibﳮ�^�?t�#@֐��1�M@�[˲����+N�9b�|���¬Y�z�0�bW��m� ���O�����!8���I�*x��w�@��9r�'�F�,�&'~
�L��CA����� O�3z���ap�� ��&�}5
����t�*��D��.���������x����	t@܈!��N������n��<�)��F��
�>SZ�~�\�Pt/�1��ƼWO��-J(d�i�;�9�(�RI(:rݰλnW�YPsbx�	���f��c`�~6��X�Ӄ�z���:��}�	a����t�4R#�8p�ߣq�ĆG��	R�y8e��;ݲX:8g��Ε��n�SSC���s�#���^���ӡ\k�q�0�J��
1��h˩N|�{�Ҍ��m�H�B�+�q�=z���eD,3�饌�!b^%n@���,�wm�r�,��&t��x��>��gd�e���<z��X��5�Z�[�(�i�G�ql��ĸ�J#f/%u�/�9Ŀ'�v;{_��0"���QV�c�e�>_�$f�w-җ���{�� ����7&�H�9,K�����	S&'��e�47M�����8d���L�S�(���R��9]��ȓ���IXuD$��\ �P�r�*�#Vl�y�6K�L-h��oOQ5��eunC��6Hió�Ց\=�����Q�b�V,��C�we��b
iB&�(\��;�	\+�F,4c�9;��W8 ������_:<t��D�����W��[�|ʂ�]o�쓪ˎ�����8�����y[m���1e�c>>s���U�\�f[Է�5q��<�_�z��[fm�-H����%�q��X�uob_6�hT�&�2�b>�&��.�������Ԫ�1+7��1��<
Jiy �C���^/�����/�?L�yʈ�e[L,y�!��u��OwB1s^~|O�#y+(n���f1�Z3���U��RCy�mc�҄A���m$�N)��~*d���ˮ���Yh��2҇�f�R�2�R��ȵ�Nc��)W���IAzБ�e��`�Z6�|�cQ�<?���A{x�Qq*@C�EH|�^H���eQXe%HZ�A ��ߌ��<���%�<��vW}�_�6j����]�2o�"�K~.&`��<��湜T�����N&;�+X�UHB�ƚe�g]�:����`����ǰ���T���(�´��'�AK�=����h�x�M����+��V�e.Efp��_��Gx*�5�Q�;w)� ���F�L���S�r�3%_2��O��4�����=(tދ��4�-8v���o���I0���W� yм��:L����$���5�{1������v�>�{Ή���j���y�ڴp����c�Ď�T$��}Jc��`�=c���3��:��W�&��Պb W�Q��CF/j9���5'd����c���0�]�{�|�Җ�M�� ٠�]��Ѥ��ėF6�W&P#��u I���C��[�x����唯K�Ƃ�"���`�+�|R�g`��t��:5����V�(��2֢��w�λ{
�S��y�_���4S	��(0`�W�����#�X�)(ga>`��Omn_s�X_İ�6�7�x��v��r �~P���Y�q˭�.��+:L3-���p�b�/��{��Э�-	����c��]J��屢�\�ߎ��ĐO����B��_d#�m]AQ�ӳ��@�B;5~J-��GK���j���Tu39 �rO2���m���.3紓⢼�D�_��k�p����)ʮ�WU�ۢ�T%�}�@��\�v�[�Y_ڰA߲z+$K5��f�#v< eƓ�$�\�����3h�o��� �g�{��^�ƃ�N9~+Vl)���p5=���-k1�h�X`h�g���`=�s8?2�o%V�S�p��v��v8z���V���O�׆qRץs9l��:����in{C�k���ȓ��ɕ�����ʣ�Im=EMQ|!�����"	��"n�u���-K��S u��XRa�@�����B�4~����oH�ҋ��P�@�ޏ�wϓ�*HZ��s
Xo���L����M,j7�M�����dļ��
kV�	��/�%T�E�^m��:��@G����4/�^f�x�v!��?��g�2�:�[N�y>�V�b�!4�d�a&��_@W�/��g2:곩����in�(e���J��t*����Cb��x�h��鶘d!H+�n)�"i�%c���Ts���&�xg�oR��$�2�����\u��;_���+l���1�<�H�6]�%�/7�)� w>�5*����%�z��(��QX��}�iB�u�Y������Ui>���:���3]^�����	�Z�3e9�TR���Â�D�`��[�:�g	���<~�����{͗��b�`���wz+Q�|�<��v��ꗙ�1x���Z�e� �q�٦0�FU]��E�qȞ����f��ݧ͹���m�^� ���6����"�X��B�}�)�q*�v w0�?�OF��HQ{ԛxX�����۬������FU���`����|�����N��X�Tr-�I���=#��Mo?/Щ�Gu���&t�J|�%�|���{��8P(t��.�� �
�m{Ip|��ʊ�aU���%W����f�'	$1'�<��K&˶4�{���T�.�vB�Xp%��L�96�ā�v����?͈��l�gC��ajSэ#H�ӽ�TU9����m,��;GNY&�6�c+)x�iW���mdŪ�Cڈ{s�$�~k����c�����#X�Ol(��|T8m�546I�~0���+��0�՜��N��i;��8z?���=@J`�e��h��^ZC�U(-�
�
��k��}Ԫ��B�<i�:R󴱇�!��-��v�5Ss�G)�����b��b��4�h�d���$5�%�@GK����;kr���z�1:��m��K'�:u�w���|��~��Ṯj3�Q��|�~�
�>����3D���Z�rd��q��u��R�
}K�H7;A�Uy0�pk�|���������T�d�ւ��YB0����O�� �><���c�A:9�f���;Ѯ�H�k�!4�ljs?�A�Ǩl���i�"f��b�
c�c��z���+���p$ߧ����~Qe.W�>�:_��&J���5�*u����Hf������F�Աi xy z?���ASL�98�~^	�i��X�����۰����)J�N�L��9�-��0i��l��Z�pݓ��}����xhqӼL�ȁ�;�[ۢ����\7�~���s�����Ѓ��#;����l2̤�j"�1��g��"�~�����+.]˄p�`\���ݒ��c�)��]Ll{1�ډ�cI$���b�m3)șl���:�}m��Bz �J�4�Qc�m����6�q"B�K{��/9nN�rV�U�?Mi��kX���mu�����k>	��ixݑB���l�8�t��K穹n ��F�ڤ��-G�?H���q��P%��n9��LN7�W3��[�� kE���e�GZ��=���j�	����_�3��<�0'��HK��wMnN���];}#���Q�o�E +'�c��^\ŀ���7�-/pJYA�w�<uΛܿQ[��K?%a�"ڑ$zP�]��7���9b뷿3kn�5t�SQ1{��%����{Ŋ"!�`�?�	 �,uiNgsVƽک��x�~wO��9�P�������G9=f�˖B�\�[� �>�k����H�!�mlK_�^�;�A�g:�G�@�y��n�00�Aܰ2���n$���
����$���p�MTW\��m�Î�e�]��q�u�%�qVS�c�77��,\�X�"$�6���8C���I���aG_����Pz2q��7��g	��j�� �ި����cJ�(���4�Q:%�07�-� �&s���'}��{�͞ިo?������b4Px:����	�ȇ8S
uz�:A�d�p�Cj���{7ٌ��.������<�J�$���o��3z ������O�<�:݌_�Mc<8�ת�z5�b���.Ĩ
� ��F�I�'8�_�,5b�u`�U�/��2¤��܆��@����ڍk�Ėa}�Ÿ� m<z+%���ަ���l�/��P�%�I��8�k�R�����ۈ+j��Ox
̤gKp��-����x��B�O��.�gn��
���{�������)�����^����$���i�oGk�|7�`zT�,��><앦q��� �\�ZW�X&�.Loݖ����.�ybi	Dښ�t�q�Hp�9��(jcD�'�2<�K�~��ol@�n {�r،�[�Kgp���aLy.oLX�]m7�(�n��V�l�F;��Lr��e� cR�O�wY_�t6�b�olQ~�b�l���A�r�w��E��	�N�y�k�l��!F��oK�a����35�s5&Ш�~�����4�r�@�}�ۑ��j���8��yU-
�il�dy�gV���gt��u�#"����0��,J7�f����Gqp���
JnEY����?޶�͝���vt��JX�Xi���>eꚴĕ�Ũ���|$c�`ai�ͪ	���%#k�����Rp�(�@|�΄*�F������/]O���_�1}G �{a�������3��;��?��[`��������X�f�(����c��K]�+a�`���n΄�wVI��'G�����X�;�}�8(~��,0�Le� �&�I���'`6F�;��Bj�E�����)�!���C����������tl���d𔸠�(��=̼�k�˝]-ˤ�j�4U���?7���r���)��4[Γ�U�8F�Z���α�/��{)���Np�+0�H]��ք���:bN�ڢU�H?�Y��}n�_�~ѭF��#BW5�e͘�G����
�]���j�{�Ƒ�T��ux9zn&B�G����*��� /\����K��-C��A�k8J��䜽}�(Y.�x�QT�a}�:.a�*��xɿD���@a��#�^Q�&WGl�� ()#`b+�[Ã�J��F�D��� L���q��'��[���G3C�k�X9T���L�w�̋��w!pd0�6R�A�/q�����@S�	1��$�۟6i�v���J
���v-~{�˄"��GӤ�Mg��sN��!"�#��o�&��@|N+N�N/=m]8��o��5'm ��(�6����ئ�X�G��l�s^�ª%��k�����*��`�KŻ��!�Vvꝵ�NH,��;���n2��W/��)�S���J��x�z��C:���9'~�T�D��ϏKR+?��Q�}֍|�A�C��߻^7�����t���2I*��X�-#u�T1s(��_?�(��ć�J�x`�A�T���C8^!�5O�'u�G�1�PZuo5�v�7J*t�Fp9j�� ���J�Б]x����z^�`��*�q`mF�ϖd3����?�����ؐv3�_9v'ϻ�M2O�EH{�IF$��շ���I�q���?���ſeICòX�cP�a��'P�Vw�|k� �A����z����a�Y��`��.��V<%uH-�ԏ����r6�˘����;p�Xgz���i�-4�-e�����u�>�G�q�՟ő�o���i~_�7H]�4�2k�F�#r�V�Q[��4�v���'���\79�.�4xD��]�����?X�ß�aW���L��x��Yf'���B4�kϴ-�|�,�U�7�=�gC��>�~f��y�H��8��p�W�:8w��aJm	���q��suo����i��o7qmAy�mn2�WW�3��8`xHk(.��q��ل�x�Z�%˓d�)��NI����ӵ���P�v�o�m&\ΖP��l~�-6@�7+ȉ��!iz�8w�7د1�{[����.k����E��]͐��J ��zDH$sib�ڂ(�i	��ݤ���&u����7�� �b�7΢��ܥ�<��m��;�h��x+��t˙��	b`=@�:ԨSU�`���_��~L�J�$�I1F�2j�Gx�j^�$�ˡ�뇍l�Pv�-��ʉ��QǞ��|4���~���!��-��w'��P�1�)�?Q?V��Ow���v�#h��U 6� S&�H\��;��-X����xff�ȊGI$��7��b�tX���_�Q5���ξpI|تQbD�;��(BSS|þ�4&���b�=�m�e�ݎ�K4�r٭Wl�#y�:ԅg7[j�� ��:~y	�a7[��`�(�(Z5���z)}�&��O��ґ|����I�d�i�+���`�ᾴ�b/Hv�_"L��0�a�ڶRK�+m�4��vƆT8YB6'�m�M�-�K���v��ĕ���0S.î%�D������+��Uj
�{�n�s�}��X�J1����q���(*���(��H<�D|��=��'5z;��e�
c�� n�p\����ugQM�fV��Rơ��EoB���x���%���N�Ӣ�k�=���Օ�R�\��t��+~`&M;O.�i��]i&�R�	�|pKy'o�OdS���\��"=��/ ��n���G3T�֪�[�!�Ї�C~p����\|ְA<1'��d��� ����f��Ӣ��:l�s�R�r���8���@�@���I�Q�zU����f��cy������7Tv�ϋ|�ةW&��:�s5���C�f�:���Z<�3i�c����`L/>�.[�Kp̺n��+uЏta���M.���YP���Okt�����ZW�h������o����jjT���,i�1����i��z�n��n�հ��sۢ2�hYl��?��J��L�[Okf>��2�7{���8F��U�d����q��y�����޳���J��۶s>/�1�ȣ��v����u�֫�����_� ���6+������oǼN, A��t�����L݃���l�O��&zʩ�2Ă��>��	�4_�3ѣ�pR�����I��Ř}����@��H��(�t�D��7�MVMc�Z,��m$�Ȏ}%?����d�w�)���Ø�HM�F
�\�v=��Ľ�t.��rX�뾳>�Bz������Zfd�����јri�L��(�?�>�KO@]�eB}�~�#�|m��CYxq��V������p�qE"���D)c�������b��R�8�W��U"r�E�HnԞ�	�`���#���N뼃��H�|�q���	VO#y�3P6n8�;t~��n1�t�P���\C~�k'��)���B������b�,͉�9S�u�g����v\��,*�!'��&(u��@봟O����TE��3�b��S���g�p�ŗ�Ay�_մ{BJT��"':�C-ka�;�i�&�����L�LN�ĥ��\7�/��B�f?�Ŋ�[�ơE[9�����CW�i������j��@��c��J�ݘ��ۋ7^�3O�����<�k3�ث?�e�%^�04gd?;�X�L�Q���1�`jG�����t�k}~0�%�d����[X�8J��@�N�C �TdO�쪾��q���������#]��^U$J�D���1�Z�p�S��yȰ�a�n#U�wl�~��e.��
Jپ��O��q�a�*!b�<����Q�	�
���&�$.�B3�ҍ�KZ3�6BcrZ�խ�UqɐT��n�;���`�����b�#z�9/�k��X@Q%;C���R�X��u�Ny|��cZ�e�ۃ�ru�kR�3�Q���sr�ci$p�o[ᛊF۹�rfT���Y�B
TG�>r��.����4�2�����-�_	��B�ۭ�-p��r�Nf�Y�ǊK��i�����q�`�f�ڜ�7�l�f��rw��nG��w1pӔ*�J.ʞ��٦��L�7S��AѳR8[��+MVo��WS��}�~Y>��=�w�8V�Z��S��0���M����` �F�@�^|�P�����nÔc��0Y�=�+p�OEA�TW�r�	1I=��t�c,%N
-����[#��K��(?p[��I7�a��ݐ�����a�`E�	�H�K��.EEF��9iu�������y�zd\�,pD���D"��~�����"$�Q�(~�%�la�"���1+�Z���]ܠ��)���V�p[�����`)gJ����	&.��Ĺ%&�YTc�95�'ED����e�_��Q�P��t�F��|_L;�(�e`�h����%r�����;�F��J��4�_N"�p��3­\�2����(�N�u��|$�>�K.sR���d�긌��,PUެޟ²����%�Z:�˷.X�`��\S�Z����/I��lͫ�IŅ��l�O�,��%7��%6a���M��vh4�ԾI�"7w'�鸼@�=�ʡ\>���:ᵉ�3Vc'9��)�s&T!6��^&��_f��H�R�W�\�6���6焃���XsJ���=��M�E�(����@�b|��&�Ut�fF5��8�T��d{pK�=��|�E�-�D����.���"�B�{�i|���j�ap@���H#M� ��h��B�w����U�ϵ+���L�U����R�*��e⤨!��i1w�]|`��fW7xv��6�
,�KD��"Ey�#�N��٧]J<�*(��Y��*�E)�A��C.W*@���kH�uk�Xy�U��Y�5N6>�sH�s�h
P��C��x�Ì�m�_(���i�ǚ�!�WP��
0@�
��2�N��Q��=�\9c�Ws
��~�Y�Ie�k�9����"%�ٰ�~6`�����ݎ>�W���w��ōn3�Pl��,E1�7��LW�o~$���F_D
�Ѡ�	�E\��ÝW��?���ݬ��B^�dr���avlNTwR�@H�#�dP�Ŗ �Md�թ��(�G3w]�x��"���������-Kѡ�ή�� �pK�úr��]�C�˞����=�� ����O�$
0��n����=M��C��jfu
9�!cٙg�D&7&$�� /�zy��,lb4L�I}�E�.��9-�D��̊M/��K9Ws#�x�E�-С��|���-����g�c�����mz�`\���i�Dw�Hŉ�]��:i�[9�ޫ���f�B��̱�����Q���x������i�)�7�=���q�e��߫{�	M�W�z��;B@����+��cl촍� |�)s-6:Q��4��%z8�!�_�`�6l��t���!J^		��r��eW׸{:)V���)ƕ��2�|���qO^�o"�'H�ٌ�N���/-M�tY�.�IP��l�7���#�J��C\�#SN�������͟g_�(ʝ���S�6��f���`�e��'�	w.�K���HD>j;�<�>�.{�N�(����*ԗ���7�Ǿ�y�$�ʀc�j�`��.�������
F��u�c��g��鶼;�2N�hvG.L���)#v���4�u=J����g��(
�O�<Q�ʘ�.z�ɱ@c6_v[�C	f"�l廖���U�'&݊J�iQ��v��p��p�����'���	�Q<�W���=���,�
Z�4�;�;«�E��?��l�	C��;��H����A+�٫}�T�9�ȗ��2�i۴��J�;�C�q���;����ׇ]}5�G�%����c|�1��Z��:�����K��nWH$?�;�U������p'O'_��A���pHɺ�U�j�z��w��6_��067S(��颧�y���X�E�|�y��w"Ӗ�VhE
� qب��	������%#;W�<y܋̏����z�WnE�%b=��3���w^st��sj�t�݇�t�W�71�(�l�Sa��&�Bt	*n�\��}t��qC�f	}����z�#�﬇'�K�L{�A��q�E)�~�
^�9��7-ǈHkAb�	/v�cx��{8I��⋜�	��t�f��&��xڵ��5,�M�[�����I���7����RHT!��:LƂl'&շ��Ma�m�Y�N;!>[]�Ջ��r�:�����8��,YZ�F}��=
��l�����`�ࢹ�(�620���l�`*fu��:�PQ�u(���xE����Dη�{��Z褱�%�S��u��_Y�f�����~�;#�H1bր����Sٍ{0���=�'v��{8��]P�Q��K��Ia���!��vZJ�.5�|Ĵv���g���;1R0��;Nm�Q�����@�Mô�'��Tss��4#�����FK�fVuu��G
�~�~�Q���th�k�� (j賣R6�C���4u���j�K���Ц1�+���f�ɛ��4��6��WւӺ��eۅ�z-���y�VjAOu�Y�uÏ+�>�oE&�Hgq�q�W����]VS��>M�C*��lkD�2\r�I�;r7M�,ʙ�@�'ܚ�r�SQ�%kX�J��O�M6�Z�R�jr��1�Z�CD��h�	���˱�H�����;��y�j�qoy��*��-֝<ى_+��0��&�h��K��S�|T����1	|2��$�z{�A��j���t��H���vZ�h���-������r�pʇ���#���]߷#�[�CC%D����D%�yc�r��#��8ie���	r��!�-��Ì9�ov&I��KG1p�?��Z��&�)����j��|�{�����B��R��K��X�iMM[�Dy�εW~�f��;@��w�j��@%��n��	t����y^J$�=sh��~��u���Йz�j�`t@{ }h���}��d���<:���`|�n�Ha��	����m�����'%ޱ/���sm��b�ע�]8G�m}�MR��j�ؕd~>�s0<�uq����e��:�>�O\Buh3�m�妍4����$J	��i��S�^��qѭ	$/�Y7�h�-Yԗ��A%�I:���k�xMy^�F.s�$�z�py�c%$ ɋ�g��9�)0�G���>����i)ً*"}���@	!�#V�D`� ��:���l}YWi��`q>?L;��4�w�a���UV6�b�tt�B�F��u(�D�Yi�`>�%�@S��]5�*i�D  EW��{�U�tԛiAVo8�0d��E�8���2daY�ɢj��fM��Ĺ�
o)������"���_��,�QE��0��Mp����L^��&���3�v����u.%���$п!�b�6��}�=���Ȃ�v�%�ء	��� ����6)�K����P�QR����ޫ��AU�4���V�:�\X#�1�$�#�Ɨh��8���`��������%+���D�9�L�K��F�m��{�*7�0S�4���]P�=�o�ʝ�D��UQ�|��p/۬�V~U�ND��v<�Ϲⶏ-*��z���S���=�ZxޗT�6�U�S�M�=N�¯r����UX<�M���ANJ��J�$T���j��m
��i��q�Yaph�4�� �0�e�-V�|�PON ��8Gh_�#?�(���1���aϟ����9�����-?|K����Q]N�aȻ[���,tl����1)��P��DԴZ��I1
���׌P�]4,y	!�S쑽�x��%��
���G7^�";$̈Ӭr�O)����UU*�%�XQ�گ� 3�7`�
j2�˿ ���Þ�Y��v�y�a�=��,G+%�O>�s�S�IIMW)xQ���������t��ҽ��Ni[.FG�fj���;)��-��0��(]������}&�Љ�<��U)}H
X�4e\���Չ��9U}|XL���!oD;�q5�K�U�	c+F�% i����K�u�zZ	��6�<�&�Ms�f����Q� Ъ�#�q~.I���'X/��M��ֹM��2(���ro���f��W�wMv�?ⓜ�V��6���JF�ᦸ�b�O(���4�L�E��BKj�q?C��X�Y�b��@�2q�6��.No3*�=,�x,/�y�7�ľ�Ј�b&��5?D�7lC�ճ���$�a/����2��^t�{�ͅ���&:78>�BZhͮ�ojW���b�ŲA�1�r�n���Ќ��8Ԋa��ށ�6/�_q��;9�0'�Ŀ p 8Y#�D兊H�f��A.1Wq��g�0����&S��@�ѐj\�^�3'�w�\6<� �MY�F�4�an	�� @��pC	��o���g��_��AG����69D:6^����@	,��R�/lf?�z9ڻ ��������z���\�b$�A�d��T�yI��a��ܮ4�<�����Q!("�C��3�u"Lo�EG%�[��C&X/����nc�&�X(@��<��@r�~�U���Yi����:�#O�@��
��!r��y�!u���E��#&����D����5���ڨs�V��V�M�� ��W)�z�I��� �!Ez����S6�5��"U�dD����+�i�2sε�=�KO�������/��):�ڔ�=�
m����B.V��n��hk�f��RZ�ܔ>�V�����^�)�1|�?�c���0��H�� .�6�yu<�Օ"����\!�*n����D̽)V�km{�_w�8��	���P@��E�"-?��>4��q_���
4	x��Q�M$w���R��-��n�h"1��l������s|�[��DY^u�ff�hFYy }��h3]c��h�"V:���Rqg:��#bݪoeV�o����w�Y�gJ݉pe��9|;g� ��%$hu�"���IT;�/ɼ%�W\�E����-\�T�Ė��8v�)S��lP���ݨ_C<�J2���DӁ)��X�����7=>�r0:P��ܲ�lq�Ţ���Q�sJi�Q���n�S�u�l�N	A,H
p�2����+9�F�K�3��C�Ӝ�w����=�~��t`l�Ɲ���5r��e��
�+W��ݱ�g� ��d���T�~0:kp��%$�{�����G
Q݂���d+�dz�՜*�pPQ�*�KB0X4i�T����:�q�ݽ[�.��p�8��#Ki�1�z3�L'��I��p!ל��;L���<DTI��W�[#[��_��́���!U�q(fh�!W�ɛ�S_��q쓵���åA o�c�o�R�'��U�,Z�}D?1�母ȏ��B�99��CQ�Ŵ9��En�;Oy�&�m��3`p��ծhoH.�A�Nv�$[ϳ�bK��o�m����0�*�Dh{�E!�Yf+*SexmM��!����^J�>�5�+�+rx1/KE)����8J5������I� �0�5�yg�ְ��.�m�j�"���<Fh[ky_�x/}�0"�o6�/�(~��}W�	���VȌd�o7G��� ���8��k *d*9�Z�����U7f��Q�p�;��>���;X�`�G��|�����&�n0�7��-�b�	d່J��x�z�L�_P���a�Ψ"�CV�1��ő�	�HG����3��v���RgA]��ꅓ|����D�/���W�V����8=�E�9�B9��}ʷ�g_߷�`���kD�B'��>Fл�HAG�
��}�\D��?EY��8���(=A^��D��/�נE�5)��g�F�o���*�Mc�5�����KJ*��Wb�;�����ul��Z���pjْ�v&�_sމ��k4�	r�+���¿~Y&ֲ'����p����a�N��k�v!�M|�c�v�ju:C�'�4H�eW	�>�cVԎcą���g�[�� �sg%����
����Dj4�OQ1W��/���c�jQ��	����ٻ�I��i�<M�D��PW�H�䝍v%=D�G��fC@��Mobљ���WCcD�D^�~*����4��l���1�-�����Q�F@��ʮS�R��T#�֫�K�عD�#������E]�&�z�4�f+��j׷@�e��q�r=�^"K}7���ʎ�3[����b;k�r��������L��6p��N����.�s�2��P�>ɜ;8y���8��_���`Zj��鈂̊ڻ���Dx���c�Ύ�l�A�QY�##7HxG��Ï[w� bj��Í��{őh���m/�[�+UY<�:�k�{b�=���e�U�O�4S�����g�I�2��+��e����� m����y�˱�}/q��⻐�I��?�'k��9��{!�z�-e��I���
^�؄�S�.VBKdPB��`>�����<
�5�&h�����q��/v�Ȭ���H/�����tOư}���:��A��HS�<��ē����6#�h������ޤ���6#E��ܻ�=�C����m�s較V5�h�[ҿ2k(=��>��F(��/L u=��>�V�2�n6���v^�=���;4�Zf1V����������+MqCQ�Z¸���f�?����L?�c��u���I���8^OҾ�F[^?ΦN�)�Ю�ǰ��q~�����*�az�`�8�F�/�ҏ� ��CC��M)���~p�é�̦|$\,�ޣ%��;�@2vA���foaXX��}��&za�Y��Lg��v
��Xe�����.R}��<}Ip�*�z��c��z����Ok�CV���e�X"�%�̻���V����������1$İ��㽖��w�W�BϮR�p:A�"�b��Xۏ�Z�$�  j��v����c�
��$``r�I�3�,���5�ݔ5�`�a��(��Z��:��o����.Hk�~�4�@f�|��?�[�hj����Jmn��3�׳�T8��� a�pm�˘}fb1D7M�2�?�i��Y��Zr'v�nƷ�<Ւ<�ڰM�"ń�e���q�m-�`8�Ճ�O��p��]�����!�z1(熟b���jb�U>T�Rj��e킮���/�@<�R�L�a�UƠ��StZ�=;Y���Dn����,`��|��G�&���!W�/�?X��RR��Թ����n��t:�M=GdSml��@�x
M$��R|���(
P�����,3�=D��,�~���6Y	���f[Z`�zE9Jz�zԕT,,�:�y���
��5w��I5z�PG����sZ#եUx�`�x���^+�z|imo��^��U��*䋂6�XsF�����6�M�{�f�7�|��`p4�Q�)�
?��'�ۮ?��ХZ�x���:���<��]Sy��D�>�"r^��"�Ċ�Ԏ�����=��)Е���h�\X������d>��S)d	�F��u�Iz��Vn�4�,��aD޵u���X?-{�k�O|�&b����&��%rG��DhL�Ϳ|�l�x_��W�=j��Յ@{�;=�x���r1���2��x��ɵǣA�R)B]	�8|!ආ�]�b��L��Ly2Խ�t���9�J�U��dʺ"�ޜ�Y�M�_�T$�!��A�J�Q8tֳ�fx�~F=KO�K+��׋X	+hn��X��}��^I'���*I7���ǡR�Nd��P��`ʑ"��f�$�$L�.e020���xt7(k����I���s�c�u��y�@�M
��-r�Ջ���4l��ٽ󬸺�N�B7'�fw�&[��{���蔫�"tO�`�ۨ��F�i���̅O���j-��ߘ��!��A�ڕ���b\�~�w��l�l�T|Y�Sz��@�1�3��W_���^��֊����hJ��.c��="W6emJ�Cu���m,� �Oe�S��p<&��P0�	����,��`X����٩�J͖;eD���K'[YQ�`�����S�9к�>�oR�Z���u�������~�H��֐�=G�HW���/��^3�'�q�q��tu�b��ȹ�w�*lq�z. ��:�H��G��E�)�9��Z)���X G0�Y������}��2i�X���b��&����8�����e�#,�^��a��kW�V���]K��4Y7��S*��Ct^��.��i���(V��T�~tgN��֌�+��ۀ��N�an8.�A�W}a� Y�.�Ėj�Vu*�Υ����TW`V�:��Xࡶ�a�-a*�ɔh`�X����T�J�����p.��p�m�.�=�/!Su�5�M掕TY�k����
��[�S�ӧn���3}��@��]�|��g�Q�l��uR�����΢�X����E1�z���� ��6��Xǡ��a��$�]C@J�L����ٳ��Ӈ�W��Y���r��l,�p)y�Ucptv�|橚O�Mhؓa`B��U۪��k�:
lxr��� �ڙ���)<�,��.��vnb���}B��5}ys�D �r�����1pr�,�m(,�:�.o	�.�[�q�3�H��~0��:��Rqj[Q��(�a��Q��
d]P���L�R��Wm�hq��V�7P9���ǁ@�yz���D��ۭ"�<����_�<�$I��@85hc8� E&S�̴�W:o����L��SRT&���n����3d1D�O���u_� �@ ���^��֓���� ��q�v���d��N�U��_�\��yÒD�S�`I���}R9�mR��g	:� ��Iٝ�Pʋ<�������!�(a��,e�X`uK�_��j9�ZǓ�b��ki�?
e��h$Ծ�N�JOjs1����<�p'v��`���x�GZR�;\�ܿ�+�
�/%��.����U���	���h�[�P����%^:G�������.��9~�S�iW�5�@����L����<���fE=xqV�H@�u�R�_�!��z�"9$�j�$x`lȧ���LT�aN&CD�G��	U�S�W�S���/�HX�O+���w�/��
x�!�~��h�?E�Ƕ/O������\�����z*����XN�<G�p��1�>�z囿RC?Q��:��өS��Iʘ)�����V� Q_��z�+�὞��v@i#g�y��: ����[��h��4��O����޼�$	-�� ��0�&��~AD*U��`^�V�E�Ŗ��&(1��	?�<��j���.��y
*�~�}����n'���dzȂ�r���G����pUȚ��~.J�"�w��_^>��V+?��	1y������A]
g/�_��W/���i'QNy���T��M��b����n._Oy�lA:ښ��&�� �QF�������Y��N�>P]x�q�G��� ��.�聒mn,�x^ҬE�R*��>��h7 wU΀�}�H�X�sLs�H�������6�tq&0L"&F�mz�O�x�x�#�Ja��S��^��Q�N�L%��*�@�	pe��׮* KTԲ���b�ixWC�/�3��6u)��@2�s�J�;�=� Ug���. |j$�&Ј8��<� @�A"nˢ�tޞ}���j�2"���/��U&2��5em���yCI���	��M��z�0h𿥈�ߦTa���Fݍ��d7nZ���`A9h�D��'޺~dM����Pg����P�q�%��6��v��Mԯ�$�U�;�0H��L~�<��յah�"�c�o��`^�ޏ�.�9�b���p�;{ɧ���7�.���ŋ=�t 2z;�4�dJ��UY���縺��S��h����z�w�>�y�nٹ`a�::Uf 53�w��W� �	/e�sf���kਚ\':UcG}�N�C��$LX�U�-pL𰚈1��W!Y%��݌�p��c���Q�&	��N0���ʬ<��3�{����$�g�I�pǗ+�RE&G:�:�Z.��Q�g��l�U���<}~d`���|��؍��� ۘ��D-�4�B,
s�	����ΰ�"'͉�w���oO���S�s��ydA�R�ѭ�|p��@��
8�l}(�m⼟B����W�g����������y��_����U�N �x�4�Um�W��0�����d^Hk���'(������wj�_�t�������i���6�A��j��R�[�(AAK �;!�Ĳ,�m<���}J��C��i���&L;f����J����68O��6���V���m�m�!g���k�0��������Wl��)ĀB�Aj���B�W�V�,!�><��.��be�
Ci��d@�8*6����x�c�9-2j�zUee��\��1���D�Q�+vJa�?�d�Y0�ߛY�����f�Ƌ8(��W�)c�^�~B��%x�MA��²�t�&ll�I�9օ�����Hȶ��G@\M2&���l:rպq�n�7�T���@`�ji�ɅB2�t�d�ʓmQ�zL��� ��M��e���������]@�d]���d��C��2��br�fE@$��Q\�t���Ъ�s�k�s���s��H'�;-�Y��V'A��-��|)�lzЯ�˧�
@4� =�>{���f�����aG؛xH���z��q���X��o �B
aY��/�yϘ�6�:8Yna`
V���c#17�E������\�C�&)4Ru�o������+�h���~�]��t6hj��l�/�a�jڰ98����Ie,������w��_�*�OCl����C?��E��|D'h	��>�x0xY�0�F�2]n;���M+gw(sct�>]5��Oރ�)1k0�(��p�n�� }/�uD>��ً��_&��Ҍ��O���� ��%WtUJ��A�_�r��"��76YT⊞��h7b*��]'p�ݾ�d�=w�K$͕`Vk䈠�ꏚ�"b�o�����C�!@H�흙
������G&M����?�2�Sn��;���o%Y������+�&$���H�yiu��4-��)Dr�����7t,6�y(m9>ʏ
���S6_���P�*�D��բX4:7*�h�ϵ�s���W�/qʦ�\˲Ej.�c�(8���hJ�'���"�`z)�@�`39&g����e�՛H�[5��]i�-��Pw��ت՛tq���V�F��w8¦�a_ߥ-t�8T^���,��>x-{��lz����;f����~���D�nYx��^�m���[��T��_,@�뽒��� ���f��#sb[�su��dr{+V�Kf��U�͹�P��C�"�e�ޥG���ݱA7�&�	��j�sN�՚By!�S3�L(�"���һ�Nq���G'��]C���3�1l��)D�oP��#3e��f��g��yF,��Ant7���~��yef�-�]ڤmW��ri���rG0���M�c��s��:�sk�'��l|������E�"���sa6���M;6E&���D��$z�YBM�ͥ@-?Io�>9��SE�`��vM;i�A# ���[�Zd0$U��B�'��� 6c�d��Q@8�'jc��n#bi���6tj���Ȕ^�	x��D���V`�W�_��>�u+�\���:.�P���A`%8��8����T��G`p����Na5� �T�.�s��m�C�e�_����$���M�y��uT��_���XG�s����-��@����žn�x�J��-
`�d�� �Rz��9�������£O�1L�@Tc���v,;ѳ	�O0nO�X���v�#���,P��x��c@�"F�j��Ut��؇ ��ًH@������F���s��S�$����ɵuh�Mr��	����'�j��;.ȉ���70'��@7�K�j�-N�<���5,�m��`��;�-�=h��`�&�fn��O4^-�~`�
��)>���t���"]q5�կ ��Ä�$K��?��Y�o����p}C~����=٠�!�9��u��;`$��Q�ս�p���wү�'�)��v��:�
���0Ź�.t�&�M�R*�� �z%D�wl~�f��̊8jT�b8�U�2E��[�/��3{�QP�@��샙��'(���Z�Av���amA~��q�۩�:���f���m�����ڨ�F�3K+�tD��N�[���K��5���:/>�Y����[� ~�G:ȣ�A�nyb'��� A%�Mيzv�'k�d��r���p��\W��	�t���`P�⎪x�S·<���`UKm�ܝ]A����=|m$���>>t�z�A[Y��:�G�v�zj%���� �g;F�h�'t �~g�m�pg�XET�K���	���u����G�VQ��GC���9j�ڋ��~�r�N��`���#Z' ��^�Z���&�����H� 'P��PG��-��e��R~��r�(�I��4-��|`��A'A�۠Z[m<���a�V���`b�|%4�������<`$��!����[��3x�J��ɛ�@8��Jz%��B�Y�S
R���;W�v�nJ�⚿�Z���0�6%�;�Ag�I��mX�j����܎"�~�K[X�+V���f����1创{�:x��%��'1M),��)�����m!�+�O?������K\[mf#\/B�l?���W��H ��TR�%o�E�	o���������>1��/�`�'��t�s3��UQ5�:ң�n��sy�~���P�`��NMx�:%���{��*m?���K�"�tz�U{�Scmyj��(�a��B2������ � �2ix��w��C��S�x�)������6��*�'��G����>Yu�셂 ��c�ȩ��T�T/�T��Ga�"�1�BgD">�G��T�k$��[���+���vZ[����(_�	�/�wB�G�h�$���h����*P2���'w�Z�lD����p�A�Ŋٞ%O����P��ݴj����3�!h�Eͭ�;&�)D��z�'���F� ��Q�M֕k-��s/���V��Oc����L�,�~�|;�1��6�d��HΎ��;m��--4�Y����	���aLϑ�3�� :ۑзq�W]6�J�	5V�='6���Ӧ�/���?l���rȧ�_u�� �m=�a}v�G*��]+g}�I@N,�<�H���`����<�!\~��4,2�	���-N����Ly1�7�⡌�T2��z��(�A'j@C����wW^�� �-�ģ���:!I�k~���7)㫟X'��+�zq+�`����Y�?�1d��mQ�0�x�u����]���1��Z	F���";&RǬ��#���6<[�s��d_����@�#���;^g��`9Z�a�u��Q��0t���.Gp�+P?	�R zF���[o�<�RR=�����C��z!���$(�7�eK��&˃�M_\wIo����@q���� �%��6��*��b��n�,�`FdF�)2�l�:L�T'�@�mR�AI�-y$y��W|���n�}MQc'Z��|}B�]3u���:D�}w��AQQ���s��E̎��\W�S���!!�٠Q�|$~jF��# ���W�����k��[�oHVsfk� r
��A��_��j6��"�r���v&�e�KK��	CM�vU�˨�-r�&�_�j�����q����=��l�
�#a�)� T� `�zp�������D�t|7�A╁m���;��Óv�^e�Co�·��5(ia�Jw�y�����mK�5ֺ�c1^�4�e�l3���^���K����(��x��ΰ}zu˪�����ה饧����B���g�����V?�It��Cq��1td#"�u܇Y�,8u'a^���/, �/���]6�iwH��ډ/i�}�ἧW����_�E���X7>o@��D�E���*�%�{�k"�,x�,|��찃�n���} �_��1|����� e¿ �	b���TNԮ�~v2"ډ��0z*��3Ѐy��Q�������s������,�.ş`�ȖB�a��bf�rϺ&��N�h�ugo�!�U�W���J�^@g����HE��RB�q"
CaY�*0Y������86�P���q�ۗ��i����M=��ӻ{_��={ް!`�b�����^xeX��MS�$�:��B�)�/S'n�	���dJ��&�Z >�pq_Q0�ul�f_ǆhy�M0r8)�2+L]���9�p}���U�ւN۝���6J'ZT�.�!c���U��^/�(b���ƍZ*҄�����)v�䣜V$�n��>4��)�|��� ��wxe`d���1����wy?	�5� L�9s	+�N�$l�BF�;^54 �g�Ү�-T�A�u����ð��4��P��o7�*q��c6~��y�+(|UE��%�&J*���F��i~����V�3(�di�K�0��C�^8�"b�=��WH�݋{m��N��.���s1�}?z��b��`�:zՒv����F��NU�=�\_׾��Vd�����AF	!����yy���z2ڢB����S��wgm���|7��Y�Iɜ�L g�9b
�+����XH'@�'4�\F�JbX�}�B3O�%1x������R�9���Y�1��C����wav�q�J>��Z�[Q^���M�A����b�LI���e�o,t�=g`��`t�c �Ɩ�%��I����71��vU�[ݑ���7L7�Y�m��J���Њ�b�W��,�u	�*#-�^k������ݯ�Lm�	a܃:ֵm��>�k��X��9YGG�j
<7].�Q���C]kz8�Pa�%���\��,���?;e���E����{76�f�/O]��Nn�7G�勩#�[���q`������z;)En����n�"�X:hX�5�������|�d��j��0u����G-;"Um�WD7 v!���VDݗ�B�Y��TGcp����Xi��w�E���Pp���f�DrE\����7��U}����Š����#9	���/�MKv�vl餚(`�)F_vr�`l�RLק� "��MR�e���P�1��ة���OH녌%cD��R�K���X\|��Z���6�:�
�}d�b�Gã��� ?��n�CP��v�"R��;��8���&�qc/�dx���}u���4�IĒ��+��XD�K�g�!��'��L�V�J�j����t\`�
�a0d���iS_mWD�0��>�#�P�9�X�a��=�J�\�k��r��
�yXP/!��}ɵ��`
&Y��%~l���r�Z�%,@�͊�?�ɷ}P�K��3m� ��3Z�Q����#�ͧ�D!���%i��Ξ�ɺ�߼+u����a��ʥ�Ę^�N�&��>o0�����~���p����	.�q3ٿ���`Fi��
S��TO�cA���:�(��9�@��}����%�C�+f���&*]�;�{Q� �p���.ح�[��X����P����'Z\�'�J9�=�?*���Q�m�vs%�3�Gh�G�qc�s3����N�VIl�n��f�?y���~�t�}k4r� ̽_���{ �~6t8�n����˙<6�^���4���]��&�HP%ޘ
B^`�gXk�?cY�#��X���yni3#���e�@�f�*xN�¶�r�t�TU��"�މ��,�P���1{G}�V�
ZDhGn�.J�"��T����h!w
|�
���\���οs�)�\��n��f��AE�9�n�'�ik^7�B��ݶ�	��h�Ck1�G�<A�#bPߚ3F�H��-@LV�Uy��M�< U@*��vt�����v����E�cpG'�_�w����Re��N@ά!��X�|F��E<�z���ڴ�r������ ��&X�c"�:�fx�a[Ln�a��9io�N;N��y0��aSW��Q���r(�����J�>��V�"�I��D*٨�.U�o�^cQ]��Q��[8'�jkH�*kmacBS�����������A0�k�
H��s�ow��O!���3?ѭ>���UM}AY���7L%��Er���3͡8�]٦?pX̀�n|�"�So�:�ۀ����rH�k/��)jr16��܂��u_� �3��Zs�F�����/�_uUr��^�#�����˦هִ�Z{��=�(�*xŻG}�+zn� T�v�BԜh+����t���fQ�z_���7p+�>5�ͺ�:i�7�.P��~��ro�_���t�A�?BdX�ό�⹰ò:Ծ�W6��(�i<_�|_:� ܶ��]�F �`�����V�aj`�>�ݠќ�@`�-�8p��*�t��IX�Ngl��)�<dr����|�c<s�~gA�BVY�����!&�߃��:��)�.�fs�8?V����ݩ���z&��ظ�&㮚4��wY�㖞lj���!"�kZE�h�c��q���m���4�P@/몘��ɼ��u�Q��,��=&]��K�LVC>5��p��M�#��ԩW�K}x���NW�J����jQˢ��������ǻ��g�#�>5u�r�4��J��`��n�1ho��<�[Rt�Uֵ7�K���Q�	-�,��*��ɴp�k��j
h���Њ�&���q0��4�!��j���Lx
O8���#~�t��Lr�j�*��{Nr^r]���ϧS���&���!'@\��0�����.�B��:��B4vَ�_v�G�i~`��Gn$zn�ˏDT���1���V���7��[���L��'6�s��Q�[��:h�� �j%_�K��4�����p+�|�t^�IcxGU8t�)hr�}pE3����7
8���O!.�p��q��c��
�#�=f�V'ޑ<��}5�5�c��ܳ!Nؒ;�z�K�
�m���_����u�E��m���+�u*�-��NM,�J�A?�\�SaDO#�y�N[���ɍ5T����Pi������)ޠISP�� ��M�a����wĦ"�π4r+6�$�[�G9��Q�'K$M�iӹ��p��'��`Y1|i|@�.�~�WG�Se(��zƄ��������׊q$��U��Sݮ|X�:���
2�[�ۏ��$�#Lp��\��8r�R[W�(�Yh�ԛ^}��1�Ҝ�|�+���2�⪬� K�܍+�s�j�,��B �BK��m#TG����#N0�@���d�=*��_C�F ����V_�lO��X�[��4���a�t��ī��HF�Al�9�]�cY����ˤ�E�[��˕&��~}�1U��M��� 9.ܧ�D���i(�HM���X�l��|�*���ӡ�ӹ�cy>* e�
�j8Mp��n�s��?�"Z���e�"��Dvߢ� �y�K�?HR�M{�X[A��	���5�5�&Ӎ|5q�y���о�n������̇�G]/C�o������.�� �����-��3\�B��輏9q��>��K��b�2�lR��c3��B��w�H%�������0^E�af���!(�Pm�X-ց����c��R�i&szt�̩ ������y��`���W]��>���9$d���Ҭl����5a#�9�G[;2K�n��9�������S�%�����I9!~n��������dFfo�J�}"�������Be Ǌ+�A�Y���T;����h&���6��3�[��Nd_�7.��m�N�g�پ����0,=w?r�\��Y��/ѩS`��i������ ����e��6��<�;���
<=�B��Y��%�eɭo/���L��a��ﮕ�Pɐ�V��)��*b�g�vZ���K>�|�n��"� F)���W�'���gIO�p��OP��N�1ͼb�H8�߂�?�y��ANŮ�\5��$~2���f 2��&���O����v�rMrtM��,G:����br�S��Ii����<�1�Z��q��['m��ݳͲ�� F;�b�v`�>Q!w��pi��ߪ�4&kn}��K�ڽ�s�Fp��掶�G��q��p�nA0�؝\��.���^]�e�P,*�2Mfv�O�� ���fPq,S����;٘�j�j�j^F���|�*�J�`B�w�k횩S,CHk�J~E��lv��2@��(�WT6�iٳ(p�E6����A�4zy�ȍ����U��#akth&Q�*��h�װ�0 �����"Knß�a.^P�,H�"��RȒ\hDvtVޛK��v����*ʙ�<*�B0�ȏ�ٰ�{l��	V��,VV������v?�O���6Z8n�cl��u�m��oi/�̊UJ�x2lܟ��aZ�?��V���t8��`�K�����:�L�.D+�@��y��(T�--�X�%��qA�)=2��DQ���)s��9�A�,��V�Ϻ�DEޞq�p�̂�>6m�GV8�Kz�(ΰA±�"�#��R�>�e.�n�.8�f�@������7�X�6��Y`[SY�e��֧�Z�k՗�cx������k�\1q3*	TKߴ�:@캏(�o�m��Nad�PZB�B�d��4��������ހy�?�v�AY�Z�������
��D�����-���rܦ��b�e��(OӭE�����ev�n��w���\+vL�q�գn�v�
��݊�܏JC�0���s����l��+_=?�P�^�l)>�3��?��q�C1�2=�� �q�h�tM�3��1�Z��q��"����4u��Z�����χ=!|%��g��y����>a*bx;�ƱN������a���ct��T����xY�G�7�MEݖ��cwC�N3Ų豳�j�	����}�>��4˚W��i����"��Hi��~�6HE��%("�o��}�8V.��e�d|�L�����p�	NGٶ�Ld�a[n�O���S-J�p奎�/v�  vs27SͿ�!rڨ�{ӥ���ة����\u���`��S��tDz���=�̼BEY�G�q�cڟ̳h������W�Yc�iMj�x�Z��SV�0�����z�A�؂�`��Hۛm1�w��$ڿ*QD�-���b����}߉%�a�2Z���z���_�`����c>��q�]�*L-0���>G�gD�z�^֡���㊥���8>�����\�?���2���g���K����X��Rc9�W ۘ�H��Z5��+1 ��5��d�cQ�8�d��r��г���s�N�z����Z6�{��E�/A@HK��~�[����l���Ь�|���bmU���1Ɏ��"�bN:m6��N��tFi��,�\�}/��@��/`k^}�rа��Ǯ���
;���;��v���F��~e��IY �p~C��P��|���~�/�t��C���u�N�U�%�{�Q��28r=���zۧ-�> ;���Ť�i�`�N��9�J{��Ld��o�E"		�y#��q�{���٦�͆߷��J;�~���u������d��������P*�]�c�h���n�����CҀ�����nq��6p>��\;������,��Cc��J�8s�RR>�.���^�Ȭ5ؿ�|jxX>���� Z#sV̄���}L���ۤp�Z�v��tH���)�h9�#s����}�]��w�bc[��
"d�(������۔�����j�OA�%J�a�j�P�Z�t�N�����o��Ԁ�U�Kr�w7l��V�*��}����>��0��܉�=��OT�P�D/d����"���
fTLE�d3N�/����%M(j�;-�(=94O�U��|@	8��?��Q�ώ32;J������t����2c7��ϻp��#`�g��~�^�M�~���*z3#�p�M�Tĥ�z~��n\1�%f��г3�랬Z�֬|� ��G���C·%Ł]��;�]�5��
M��m9�]U�&�Ǝ7�,�� ��2�VK�����F��c�f�����A�ˠ>� m/4�b$=��?p�_�}y�p�E�T�;M�ݠ��E�F5&�`����{)����