// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A8GgI94DgLZXBTXEljGO/gOThjvVOuOUbbF7/ONHBu75AvDYpo5K9WhCu2ksZONr
D5Ho9R6mm4prSlK/qnIpebWWIfMZB5JmNj7aP9Ntl29S0miA+IHQbny4F3AcM+8/
a2rjIW1mBALrUTWrspQkp2xJSoRClxDHnsLdG+8e6DY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21648)
mJEA2s9YX+99J1ZkXJNk+AOBeGx3tW2YDu+eZuwPPndly0jA9dOil2fwG80PZSX/
0VEPn5SMTNGXwSnu/MKgljogVhQJBmuYiJW3SYcHpqU+D+Mvf62yEMn81Gehgzw5
fJEUm3cSe8Tr8LXdOcWpfBFeka0YKtDBoYChN8WmdNTZY9wFgWE3Xqrs13l4J4cl
Q/2AdtIATpDLKhixyI096/sCUKf7mlnMmS4pEMu1LXOtYLaoFYDqizjZBzRUGE7J
+y5DuHCAEdUuvAxvmTodXyScK3ugIsx81baA7scTyyD2NyGQEO0v6uelUAwPsCU1
6mYYf/gz1WUCtOWgYorfcBo9IolFFzKlGsOcThwg1WooXC/YpNjcdVW2lfg2HMxf
v3OkBNAqKkxx+BEt6NQKcCBzq+jzle5H/vweprXvSnZUCD0HAprcFgeCHkT+9RaO
ks9AOnEoIpBu8lGWVzhLpXOgVPeHR28PvIz3laWWFrVXWd4Qd+vPSI/ugg3MkyHQ
QE8fVrxY8K4nwGfdmRi9OfjHEmabRL1aneQJh6tXfEA0peIG0YpnT7EB96+N301Y
3zLqz0IP4TVPQJiUYAHZrDvHOqbgqZafqtg3cyjWX0YHWravCdDjKqG9z1xbblbT
u540nUmJpNlr4GEc2IAQqfJbVtRUYa8n8pztQvKx6wfHCFvpI4npcopR45xLKFEd
8gKfLQR8wGVfeXBRgFmK6RgMDMcBoErYmavHGf5cjN98ckkB7Cieu8da/NVBewtQ
Q8bHvZPDbGo5s1V9cpmQib3ZMnQ/FBPElv9Jc2wcYGII4QXvD5HW18wtXQO6UtM+
S1fTsl10c+mBhnF5+rIH4CxD0lP5YprSyjHhSwbUgfz7M5YZRLOn3ObRt1+nQHfe
sFIj91e7eAIA+jsCaHaLFr/q6/lqT7iBc9961DWilgj+1V/mJSZrPR/Ut30CDMf5
sF7LvCmtxJsDCi40fBh7LCYL9W1a91Xs4SGZeEOzf1kvG5Vx0a2MjwNTIGm8uEGd
FT8BcbjEWaUWpBMu/d0chaBKkemSRCcsbbcsQEj3zRjjJIny4RXarqrShqmf90QI
BoYAcAPXfpp/8ybwel6UNDfPhYXPqcINi5fSpm8QIOfoSkRQOmDAJtU9/sjTI+oZ
3NWfk8dEf4iIME0bdO7oc+IZERC4ABo8+Nn4G3YZKJndHBaMPiDVJftATCZb7UIi
PdMia9ut/8s9SGPghAuulrfG0IRTsdp3Z+2JhxJThNYQN4RZ+GK04Wcc1bjOq+tZ
cpyHQ4Xe8T9AyQ1lVb3pTvu3k6eoZ1SyRv7QJ5vF7OIV3RfQSlZsT3mnmuc3cBdt
8xqotnLZu+NLPv/H6LsPayISDxbnSrTUSPijiESVj7GzvEh9+srlDO74IU/Z1jei
p7YL0veuOsiN60EDJ5OZGBo4eeF9gqhy1K0x/0XTSy9TGmaiWR17BQYSC6Ogl1AT
lnAcKDzAi7MfHz55zWrrnDXkKm+0zFUHl9jTZJV7pcPRkzoGILyM+VE+X0VuLEu/
U4R9E45bHLXInfgwmjIsx6A6irO2JT6y3LYzZMqWAG45JxqC+iIZZtylGHFYI8qv
zZjWGxA9mAiH0wYwscNq4SD6V00dRq9QUDPlhUbz0Cps53CRyW38uRil9LHEO8K/
+NeJYZSQIDuJjgQbhH8ypFlywlT6F3Lnb6dhWDWFcKeBqZuMqwa8h/I+6FwhJPEC
sMXO7PReWGkcOEgfRQjUVKx3qcY7nzqVzfhvFrqG3vM73OgVW25LAAxfJ0rVFxCr
WiSVWNuDBsU3+LK/3+tfdAmWvmNOCrORkfMNf2DapI+KpWLh13ZwpjEgtAk6b4mo
dT9myomwN8x3BdeK76G70Rn5FX4cVLx7Whe547stko2ERp7t9wxlIgAYYBDPl+sa
OOSLvHthi0Q/jQSlCjpr0GmtCsBfdE5oUXvtc6j9ldZD9BZzLA6FfiSIvGwUVRjl
jwBb7pxW8mGvqn9IOKB8kK6GNJj/49/tXo3oACZtG10W2WWG4B3AVCmGhTtw3QPr
ZBQbd+dYuBubo2ShEj6djd8E5BZ2B8A/BdBNMdrLPm1sVWnSDwvdoKfL1LjFLr/u
oTSZBMxCu5NTzhDErPA0ojxOHTmRwsEAHg7rSpJdV+NaDLz0A06WJHM3Xav8PL7r
s62PQhnjg9z9P6k7S6cQntTaRhWkYuua5VPlRLkXGVtkvdLiIa4+1FybRkQ76rBq
se269uMh6knVuyIrC2rwQzvuedm6l0DyRU6JMyiVzZJ4AgOZ19JZVC4txrE6xRHA
vHhfEawRGYsZkCRiI1EZ4TF9NmU4DcU+ba4MoN8Ou+tzVuswzF6NooigaZpEJVeD
wnFasCrGY4Blljd1r4UHQ8XFgEryb2EKC9ebk8GLvCQxv6yod4JkJpWxdTwccXg7
tBJ7PcMoWi7wLw4PQ56odGKLNTVDHCtWLTo6DutiYWhoQoxWtVtNA4abylFnVxlY
J2724fPwUBGnTqjf/ClSw6rHaD0UsSOYIUlj6bKK10tu1Ycl9mPHW4X8UUEkG++p
Qe9tWdzWWrEc4ixEt0pcsX1UKGCuCuxjO0Wq/kTlHF+YfjJF3MdWsDl7wD4eUNk+
sZPra8yZ2wAUgb8W14FWpEpnVxanicq7MbifQqJDstW1nUmZoaki8gLgWH8xSt5L
NPae+/u2lKmKTst28GfcNpSK4JlgXQ/4+608J0y5vy94qY46Ju4Awc4bwXqNT9lA
2yC+c8xx1ME5pgkBPU5ci7oCEKr/sR5dUqR2uyOGGTspwkwl8kJjLSlUMTsjLHMW
yZ9rv1zNsA/zxkKQ7orE4k8g7VuDadYb1E74ZNeRTBj8VP1PSCKM3uO82S95qO+R
72EZehKgugrH7CUh4SY88FE63q7M4XmoUJzsZyvSb5GEY+Gku5jH0YJUmU4mtX+i
qcldsXWlTNXTQkcdfl58FPoGO76tE+W0hG7N4mvKHBcykEc60qj6bCBs8qul8ioq
e41SlAJNCNuv04lE4Ff+YgPUyv7tXJE8rmiIsxmlmlCcrG5+RnIh+YrUVHdbIwgI
zESZUlYne0tDJD3Oihzfpg4oyX7I4hViltjZIqfM2WwC5t7Jj0StqOfiFwxz10iS
EAlSJgNMcVV8wOnqyaoPFzRxsp14dMzlf8QZaS5PZe2iKfxj7C9ImpmAPBgrnJ0j
mqtZW5k5yEngGxOPS7yX8Qq3C4IQwlSAxALRWditrv/rWHDuMaDyLtxySe2QfhRB
ykMdBLayIRNI5tdwETxD26rMoTN3s2lZdXQaObaqOU0xo1F4HYw/M1q4IbThsS4R
UbptJY0j9Ryr6iQ+o0Mxu3N1ft4aNFA6awTM4fPAWf/Id2CUfyoe+KFciniNIKbw
ZQel0nciVDQ0A9ZJc1itsSkWguiNVb35JGJU1n9zDjna7bozNOfOTpLfgF9juUfY
ZWxtIX3mhwQ5d0HfuKtF92+MZYFi36P0hkPjcRWdRvaif4jdowo/4Gbs34Fpu6+F
osNqB983y3fJf0zdhb3CyNENlK8d6hrFM/eVDSkJAeqIUMxoRlBCY+XN10wqGyrX
gPEM+hvRyZCuUSI2NBxpPV7Di++VpeA9H8Q0lzjQeP1hxcG0TVcYHgpDhgfLCAbA
5Iu99K85i2wR676Wb10YBYD5xctcdDXbq/jk7N8Optv4cPKyUAQ8D1bItNIl4M1a
MVq9HHtZx+wRPus4tmUoD3f9m3mMqU5uyfCks21y7WD2U661EPX4ZRBIC4nZmlPr
jRQBhmmx5LXp3hr7BLPV44mJE2VV8Moh/lR+ld8NyiBnRWGJniba74SLuMYipyS2
Z0IK8N8nYKE1kobcn5xMneWVx3HQil1AuVrc+h1vdoWHEi2Mopes++6+61D1O05R
bXVUKenPjJGXFSDFHyqoGOb/noeQnJe+WEaILV3jdGjd0jbQZQAaA3gHOZUGRcO3
o3pi0w2gYD/Sal4u8/3yCAW5/9Leszposi0AdN98C1t8rIv+LfC7jTsrrNcWPjis
crg4//IEqwkoMo0bf1j4X9zfICUxkPQaSYqIwlPCj5m8L7+VoSLtSequq0a0ZEzK
7ytIYKFYs0WifAF8RqnnYOHt9x+lC2+v01s6zpHMs99a7HyVLlYy+h+fC9LkEZ4h
NvWAuDUp6rVkifranFFeFmCO7Spgpb87XyYtJskUDYKL8ZPh78/i6YzAe9vRY/hs
QQzYQ7q4m1VBcGXJlkIv4AmcgTUVxt7YsksWNCK3ITxlhOecbgdpPICuhtiNjV2h
5GNXTHeNsxfBDNIddZtPDNaqKwZiZJGWfryAwcsBxvNiwiUsiMdxdDEEVVWlSxCt
vkGK3P9jPnhJ/MEtPOHzSMAxM9kKMb8urp4dHv0p5DmsVeiDxLXEZ7RdtCFQDoIg
oKMjwJ3qUgeg67BZV6cy2o2aD2lsVxZ9Z82xaZaAhEEISrtRNzgitwF+lqECM21Z
XKmh4NM7wZYaAjNtkfjt/vCyHCbFKi+l0GdEY0vWl7n6CPp5LLoTdeYanjSjMQKg
whqq7XE0UmaXHSRWi7r2GS8fwWhjujjUj8M8SJGu4sGLRAxDu9+hql2fXm5Xbmib
vf+5k4pCJF8E6GqQ3mzRxoKzz6AYXx3Cx3tLFrxtMDy76KHOM+13SBL7zOrS9GrO
0Q7aoKsYuGnKZ0BRTeHowfSF+SJ9Fps6Z+s7J4Bipy+vwKrKzNoxLOSeRk5d0t+X
Mp+kzDfhtDp34ZfRQiQzTsNv57PwQcWmIE8GPvUHAVrtGw7eaYiqse6ntmJ4wRqt
/XhOlqVZ5COuerwfHZYm0fHi5VaV/WrMNiZT99Ry2qGWrUqsAvCqj+YcUGjX8gF8
eDvRDWmW/4kq9tLXSe9k0IsQqHnD2DW4AXCiMwdT3fDapUzO9oJ930xNFhU0MJrQ
1Ym6Q/S7rIUFGzC0L5FdbO9mjt2bk3ixJAnkpnoXIoPIVae7WS5/iCmMvzfT2vsb
QaIuYgCbtlGPSMBVJGoaXeyzMkngh9W+C7eDgg/D32F+qp7sGxsLPeCdUAciJQJo
iXNNTWcbh35T+5+fYunMUXf5mbw1I6VcR04mcuTjZaIBLWW9ymnvj5btjxBHOebd
iU9FzBtDwi8Fk86y7nakshNdKwS+yon4VMXalsJqN2hfBT3d0Xm6nwmbz5nVDZ6K
Du0YAkLbI4XwAAdBUU7DpfeUmQGL8cCUYMydYKDup0dFcHnCDp1nenpPp9jsZz7j
KZj8ruPgkHyWBpczuiD+MpC6pHtFV/ulhQ8skPCjptiNJpDo7mGJX5dDLBPuCglV
H1LIG6mBDJUf5Ox2begb0GPBCUFKWlhlImiL7Uy3nclhVxNRQduD5Etz5B88N3/R
sZs832P3WF8FnUP5sMk7IidKphz2ZL1GlvpKfOBFu0kQTHCS2IRPkRDuHzxOi99d
f/tGJSRMJMwYUKEPsVJFcFggIcLk5H6vwcSD/BhKFbp3K99Q1ASy7ZeaZ2wyzIaq
83tLJDzz04I7nl06rAzNy6HoIplPtkr0L52MvBIc1W3prp5eWXi5GaRfBeaNpmN3
NaFXH35PYqFxbMMQaLTM9C4OBlYiocS3eTF6DKvC26u19dDXfpZ9AwWPWi3X7my5
Xsoo64klQgTmY+ASMpZI0Oo+lax5wSyYq6IGuVDwM+foCf60TkGRSJ/PWKTG0wcg
5h09BdvtHuf0/lW3/8ae+rGcSR3Yer/1XXKeP8V0RLkkGX0b9Lj/R8t2BdPBoSYg
KAnIohsEJT/gpf8398mzAyBgM2si1foiJEjMRJ0ty4uin6HGDtpVZYOU+wWJ809S
dzm/ys0p274qnrPq4yNIpyABwmtI+snC8PW+jCKbcFDeOIZjj8dd+AJ8MfzdsuQn
C81JIPX02mBfRnEKAAmBAbQDEqGbQFENHflDcB7gXBIob7xDrEliQ0D6KaRNA7o3
1laZ3izP/O9IpWeV+t0rgYUyTE8oKMpL3KW8ytPyHcqyrV65hdCqZ+ZRx0qZbqUP
9/mer/lcFfIs3LneEjAHfqrIMOj65M53+qeita5m73HW9D1BGzajSDUd0on8DK6M
x9wXmEhWpqm7UKNU6wXrZSa9byus5pFBw7XD+QG6Z8YY2Ml8LMZAahBemc5+0F6e
2NAkNck+SZKW0aWAriwB40jLtfLntGNrNqXO89OBAd+Af5YJ3G3/chGvyDTRW1mh
fSgxsSYbVf4uRzHnPVVIEx62thdr3DZip1iJK54d7RjsoU0RDLtLhQxsqzUF076d
XwhDjGIiTiP9WECc/XuqNCBKvPo/2Yf+y5UrAIgGAWrT9uQ+WHR4CSeNfeLCJQvh
Wi4lbJj/YMixlyv+6bDUVq9MLVcDYo+/kKhtjG5VEsv97EEZPXMbQXcQTfeMgyNl
DwL1YHRyTrUZtUVQdXSSG4a6yZz9eL4OSUhQ4AhFv6NlQJLnuh4lp5rpidUOMjyX
qSWDFQ0EUbLx7mxRNrY3Cz8Ki2Uw8EDiGNq3WLeEsj5fmjkCDUQZzZD9kDdR07nM
j/pRDbxrBF2nGJMAsLVWjUyybr83/BzeP/XTYAdB8DO3n1Cd6GxE3juc6yVO3/uT
EahiF3acDMYXvyadP4wtfy6G3rOA89Rd6hasKf7wbXUGDzi8YratsRXZt9mFZLnm
S6DVv/fN1Id/VzApTeT/TdSK6SxcQB8BNq1EwziPZ1EuSj3OrKBqN4NQf/CvWIQE
4LGQ8klxXfcBzQZGzgGXVs7tm0+Rz8TDkc5YZsWHXAqL9fY7y1PrvqPdXvSGajGZ
6Y9He5+xzvmjbWrWQIeNHTVptNTbUltweojytIYn+KbGhubjqOvc9/i9UlRPBQJU
Cu0+XiBisI0lAFxsXOVxwExctow64nnEhF7B5At43f0HdhZdZF7sJQ5aDdZTys3X
F9yqcNL+OeLQrCFL0e3fqvkSx82oElC+gyCwqxE5BTX3c0B5JuNlG0rjaZlsCj7u
EA8s7hCbQx/IWeaARzkuMmPNA70AktJZamDyVvUZKjgScmUu1E+Payl1VSDbgw4j
fGByd2e5WwXkv46fgYOWbmodRZykcdFBZk9ObhO5UCbTNR2vqErU/fueubawjMXN
3GfpQ4wJJghfdCqreUejdjBt6LS9nfO5w91F0K/obC0aQFiwgY9PJOUPVjspnKLX
QmqD04O8ynjFuUF9o3fk8dkX/VfehEq8hHvFGtAqWieFWiE6t0ylBK78TyxdFKRk
raAYUIOaTTnjzhyPF3jECE0ndNjPPLcZVkuOeky7vY9znZ1Q+eBnhl7t5LfeXs1N
akL14irBWMr0DnlNHDLaM03yeP1HqT3yQaELrOgC0bUSJ04TmANMQI2jo+BPD1pj
k9iJw6oDdpI37xLAibDC7GseZ4IFobcwqfek8d/6Dpe3vdV7I/ZNGhWULV0uiwJj
GibzMAw0a/lea1X0ucadTecN8tsnsE5euZ87rly2Ou5GK9kOaEWurQwqdRnhby38
HRL35Z6LpVePth+5naepddkK2v4V9K6CIG2VNsREW8/kllgzAS1nkYIwFgkqY9eu
cGvtUi0i1CqLn424EnPJg0+tJpSPeCw4F46i2INWKM+eVoXTfFeSd7icKDTBN7Ur
DMm34+/TxAU/JFh2hQX/XoWIRD6E6aPi4OV0AXd5WXhY2qtInz0AwW5dKZJsq/Pd
maNuGf4vubk48Xmr5JwwORAN4vXe+m+EvSLwIKZbyGInaQIJRvkCLxysUV9gFrV6
JVDfvQv37AjwUSFjozKB1K90XYzyPG0TrDc1roSpetxL5ZrDt3bCqUbj9cE2gu7G
cqIQ08/Qmkh+hws5k4IWvNp6erqNpZR3/lC3Rlm92vYSXAR7AgQ/6QAnV5t39El+
tPXvFnmQtp8KsDl5T/hphWJE5fpABeS1l21WKxqlQaI4E8Mx8NNwUvxgeuDU5ca4
rOeWc6FrQ4G0c9MhkWimmjXFSNq52YnXHlXOIYXJZvMix4gRLfM2MY8xa3KFzXd3
Oh39cfEuqNtKJ4bpC8LpaDj/qXKYLXcVk7kwljNzb2CcLRpDdEDwaHD5y0641pGg
QMTVSA0FQ0KLAk85Zq8HY5y49stK2UWRYaGuW4xFPfIuNHBWjwD0wJk1yanc9wHo
+49lQ/RSEzZpy0GTjGNOlTSZXjlIAcijTCWP9qgxYy6l8Qd1evJPUSOrhcQr4zXc
SyzHrJ84+ZOn4mA/AX48d//OJn+ELPvFIyDyviHHCPO0Xzw5L9Z7Fv8iYftXAdmu
kAQuNMG2/tLVo9KdGpEEAEt02j7afXcCl1R68axccZWxV4XP3tsfKAOi5QM0ZXxa
jKKaYH1R97KtDvhlwnGkYz1Itm5edNNFZ9E8cWNhxCO0/MK+lgqgU7bFC/0Tyif6
p0T0XHNecxGKxDBSpcfQ2uCi3DjWm1sntrsSxYt0GfUTCnJv4Rc+w979VySf5Pim
yBiiYmVtkm3myhf03GeiAxs7pfecA5zJCMnU1GfzVb26aDJcBOJ6xniHjlKxXDQf
9QLM/k5dy5gR2RXkPztBkM3OQFAJKY1kafCFFmSA41tu5LpOPccElyux7bWY2aiy
V5NIMxoeyWa2n+kJlVzWIMrjEmBGM/7HhiYvfFNmEyneOwDr2Jg60Dui3rBSbW+S
jXZVhpJEHfHoo4WKpmb3yxN0g1xA5fK+IZc99NCgei3duvmTjUtSBwB7ypdeEaex
TDBlzk3AqfA3vFcDmvZVsvNIfq8H9zzubPGUA3RzDRYvEZORAhMp8tvsMqFl9VB3
qMLQLJJqlFQKHnCKqRh+chee+UOpgxrCaiBcH4RE5O9vqjYp8hiWVVCukjUMDiIO
7+O1J1QaIgr0e2gSod0s0So8kytz/mv87UsG4nVZ1g3qRCtwmFQJxWCX+hWpppvl
Jp9jPf/K/hfLSQ2rc8Zhwz5/UiifHE8qTD09zhb9y9StGQYxnj2ue0E+Y5qiAyXT
Vel8csFvsMmwGtf8rJadwuRcDXzF6X0FEBTksYOuQ66jZ7VwMDS5OQ9qWSFyybBT
Qftv8VcXnpUwPjPSq2FPq2je8T8YMpEyRGi15XdJjYRwKZHFkDHwe5uDvw8Y5AgB
XtrlglcGAX+7Cr/AKqPI16li7itCbowRspkyFBeiU37dh175v/tUr1Ld46NVMsqk
uvJgDfEJ1eeKablYVl4jAVMRQ2VTQkPqsrtVK/CiS1PODNvQdQwZlENuFhE0+cB6
iilBSuP8PiE+Nw5Wt7yAbl75gU4SzyPzPO5k8qaB9Gyo9gEXxjt+IrHuEr+vqr4L
c/4N+rM+IIzDeswXUE+LP6PqvyrAWSBcnxGN1rMN1xB3oxaglGsntFfNNp5pAqSE
+k0215gAbqTl1AAu6BuskZslbCBvfy3+2oQ1h9crPkDXWT85mgO0AX4UjdHrw5DH
e6ZMU0Vcau6/3a7SqqNAHdhoi9VQUGd4OGN6udVKYicmd4sjI1gUYXcvACsLfAT/
MxKcXglQQBE9eV/fnAW7GLRH3YuhocthQB5r0EsoapzKHhBICY6j403wazGk1UCP
RFI14o1fWzp8RgDdB7Ne7+5JU1kXi4AUyoUSS/Jc7aJIMIG+yuIPG30V9y9VsG5l
EkEMiWTmNgWLUiaX8B+vZQ9Vx3U8V2le8/K8lnij/E/sO8cyOc549Sp2cw2/RujK
Ttc170J3zW3erC/eXQAbfgiwnECo85WGAlhZtmXgrVs6ZeZwImF8ATRyGrUlnEwz
gwfe+ZedI8NTRgLPTmwVswka9SsyrVRrPAHiJS4Za8s9sOTyilCotTVSw/7YmDT2
2c0uQT6fG4y790h+yf/w9fHRzxQnu9+TukmtqUQvMfEGrppUnTT2d0Q3TpKHtzrR
IEfxlusGXuhVxXpQlY8tvgezVJW8WuZ6OCexsdyX4+U+qE8vRMna8fJlhQK3vltL
gtyBBoaK7qa+HSqFP3G2uLs2hXkBnklcVAhox7RDQhz5jWnJnxXyXHirC6jEBC3D
zI036rrF5umHMY6htZHwlG6v35C5yCLSGNPfmJPkl9OwZ/zAzxZQDBRwjvRHllES
2etfNgfv0aeSdSbbrVxK51WIo2NbVvmlh536N4BphWgeVuo4EtktVL6Dg9mV3Lr8
obYFBg/i6Klq9ACfAcEw3ik3zxNaHjmNa83FKNe1AbHFx56j/D9YafHYE7UoxxYk
To2LpH+OO47EMJK1JERDx4Xj1xGcbk7vYRMPTsb1gTufVzA/Curqhz8rvm2dOHxC
HxO8j0W4EnhFJL3GByWRMqhjqIzf8EHXE4TD36XiLnFoJpol4ro9V959qS5faaNo
/3FPys3SY+w5/T1DvY3zeeoIDVRHy/umKSXrrAEKEaULqcb/iZXpUsj5jM2hcKo2
Q4HG7mXvUexpgsIvdzLUS7Znu0mIvn/GJzVsmOFfDQNpyq/oRk7axXA3FO3BAvN4
A/nCPBcmhukl+ixejOzAJ2VgUURtv9umjqkB3sWwFZRePMcS3jsyux44HPAlN7C9
jimID2sUAo2VEhW0WCK+ry1Hi8SFe3Zfca/qVcjdmapmSdMpBd4iJTtqDH1XWuPQ
eqaz++eM2mDbLt+BLdGC9S/RiB4Yf79fh5MI7PcGekyNZmFavXnCZIIIxij6ZFcf
VGE1SI3pHKh7RJ9krdAZwwhpKUpQHMHOHka7C+k3bY9k7PZ9HOK3mZPE2NlrFmlr
yHeWLVGBf+cd6e+QXu/pIw7U4yGrSfKyr8GmrXt7vMIOqBU2YmH4GmsDBxt5Ni1D
ezvpdcLs3THg/eZSAhL6UY6Ecj3WUUmDqCGZdUX8YGB9QwGEHqnvMkLCczyg3LDf
8l6QujEk7kr6bhvT/W+oPz5Fl+O1nCTrrLVzsjwzaaIr9vOARdYVsECA4lC7BQRy
L1lmi2cDpxw0aS7+KA8LrA8iaLtcoB7lDeL3FN4qKrPxujtiyNxFomCooJUdw3oj
WF0of7c06H6OMPE2VJBTlck4mZshuBNTfU40GKQUw0/eqsGhq0NiBnSRLu2kfX/z
kVSfUdVQjI+C59tG/auUGp3s2kvn2ikCE91MJjgtNNe+3zRdhjL+iX4TjJ6qM7Yk
ltaZNCuwqoOtBYtfQNfZdqgk4vuLa3LUYUNZGl1yJYKXn9ZQDFVX8BJqnfp4tLcO
BL3B4zFs3TrhRDu/Mhl10LDjEdTmKY1giWmNy8h5oRgLMQPr7s9erws5aNZ9/GD6
8pdZFfSCr61RiE2dWXmFpECTtzVd4992555lUQY+UUaOOyVyp4xKpOAdPsJxTKmU
hypWNHw63HzpjS/IW3cEXJ3nTIRxa5uQbD9ZEGjvVYgepOG/b3DzqcfMKVVMraR/
Ev2Utq7/r0Ewesmfs7Ww/75RRKuiZIBORdTJc++o7EgqmrMI8GesjepHnwnX/6/T
334Er6mlEbXN6NeG8PFhg7hbOB0HLq+U3vbOJq1qFzcXSLq/GvL5clZbeeHbZ1zx
JQzbq7OqddrHXQso6CnMTllDcABBhJcUZqjOpDetu1pFNp5p6M+Ggo1l1dZYO2dt
h7zIipfVQYcPZze0SzenC3sRs6RNRYvjzXRntTwgVk66RHrYI4I+Rb8Va+vlINkG
NqDhvc+cOe6K2j3zM6VYXk8M2sq8lBi2v7+v3UfK6MRB8aUUIrTxri5yvpZoAAnu
QFfUeY9W7q5DIZ/gkp6omltLzVlG+dbBxn4pfQ/iRYEXy4mPSSwQpt+qRfw7frt/
SQvdy0YtBd012MsusUydw+K9ZcIiy394lKlgVllw7KqbdJ+zWqX0VgvwoJm7dxTN
azFlSFYDmC6VSE0x4m99Aenf4MZH2k9CgDRF6mzmdkH0UwbfqW4GOtfpIwixjBkZ
oYmeQvyc3EUbRn/skgkfHNcBcKe/Y471fix38BeN1azNSRlM1t6FGiXuEzHMBZ0H
ogODzuypSmlGW5t7igUHYfjZnhCFKupBiIdux/YfuMkH2PlJbaM7Z38Kt4dNSqwp
rULwPQevYlcOB3DLCSTKPU/47+sXjUTqHR6BGAPrFEXMfOLzbkYnm/Uz6JZrDibV
zmyOxecYry1oDfZn1mFB6r2chlgk6qS0TG/d6LUyMfbuhdfLEyxBxDNdoiPeNZAX
Vj1r2wq4EBGdrsAVr+qVoEuIQzz6C20BcYtxkLrwxOb1y17ZwgUV/XRglQyIfgVX
DnTAy6FghYGARbiLn7uACtlnAOoeHRJ3/wJE5BXW6x2XoyVe1zNQCQZVDRwEMLgk
bKx+42OCoOM3SHyiIq5kS+cmDXqnMDeQgomf8JddsAI915IxdQ45r5a0GLkQg9bF
Q5Gvxsqi1PmFH+3t1XkxADf+AGGq+e3Mj2jw3zbqfBPlBeateOzPkSqWi6s/p9Rr
V5/GbQynei72X9Mojozq7K+LONvjGmk4mZHNh196YowgRO3RXi/UovgWKWG1LIka
3PA8iYl+6DqYgP/Lac9TK2ybNrFCcjXybLmbiFqdjo1NHJug4p7tzvIXbnhhfbxB
QMHrjY4suynJhn23B/D8e9q9LtQyOHMCXhI3ClJvPyscrM4XxbyC13rSdAZN6mCC
QRKKFs7CPUTeD6VX0ik2uRNu/090l01z6hstVHTjAYrY4xIDSlV04luSuLHAd/M+
WTgK0iOENZaErgStlkazeixTLyZwupP0BwA1GHA3IxoCRN1SSiBVd3M5BycFrYkW
5g/66EW9rKrRKs5pFIbfh3C3P6sdgQ4D8K8GnF0FpKP2+Ahe6/3n+NcR6IHEkrHO
IqgWQBxEA+VRBfGtn5XQdIpK95MAZ6PLt7SlJU0h1oA3mY8uvEKgKjXylp61L56N
oPfr0Z4+IPxZZ6npWZbOarZlu3FiaoJ7W+vybHq6VnJ2HNMfJ8WD4p8+KdToH4RV
kAle69gvMQzGHgD0ONdB2fbp4cCio4i5hjfy7OLFvcujT1fyRo5NuWSxhpgsFSSf
dX9voVQa8CeY84dA4Z+7ozLUthXu/bJrWeqt/XTqeNwRYYM0HWqrf0ekksXm6R2w
3VSWYt+ngoekPmP3nlybSXI54bwDGz/yioxrNK6UYwjl7VAWlxX9vHOwCRkkiBCY
IU9tCncBkL2N/QZXzjzPcOhQC9oXWVWscowy0m04NKzWn0awl3xfluEI3p7v2d9z
Dded6/9+3Zpmc/h87nU757fjT/IfUS9IAIbQAORbkQAhE0fX9JV2Fwn1DCaMcS84
AIdp/58yOjcUeSo6ED3AM/gayZPQ+wTY4ujNnxF0D0F498s6/MVVdZbWonjnzheT
Lk9+vEh/5pifN7OwSQVCxbNfpRtCwIM9FQTFaDRg3aQuCXnRQsuXeQgZ49CM7vgG
9smAKX8JiOgzaCKcVKMt/14m+SIkmsgNH748WXpVnJTpnW+EzrxJagP4WSirpoZR
Fno8I1QeCZagtG10+QhklUdbk+AeOtTylF1YmWuDLEy9hgQWcSNHo61ihZ3tFpl6
hJQqBPEVCUEQE6LmVHZlRUgWvmYANurPaWtEcjPaE4Ixy0oykafExOhc3VMVYdnV
J5C+ji4GYKj2AZrokuCR5+3HmiZsTyFvGbyoL/keeUzbQsmtPc5BSYppnHM4p4Ak
S/HQvaACKyR7TcbpOUhKIPRjB5pi4NwO4ItkarDF6+r8O6n2MRl8xpnhCuBhNgFe
Tl12SuPXFruPFVVbi++BnhE/lEe1iOgmPHejDWbVPvOZVf6DuoesE3Q6KdOFHdnM
FB7QRhnPRgwec5gjL1C0OBIKYPRld/Fq9VHx61MuKfZaubq4Y0D9gvmwuqztQzT4
12lLTUOGmhcRJvzXbF8melmx61T6h3id8tDvrWINU015RXa8NoPuHYJBfrSfzPYg
2OJrKczzOdzhPRLbUmc99eqYxjga6FMT8LgtYfEZgcKbggbvWZDPNLtILsoI67LV
ht/Lps2uw0GaCbX2l2BpwX7gdhKOVYIb4JMJgtGnd0g2Rg21O111i4khHXWR6d1r
fHVqW0xQXpoDjsytcLnAlJ/Ji027Sa2qgvUkqP5IkTHZOAdhBcB2mARQwkJcBPgE
iiYv6y35zgmMX+92RAe8nWWZ3J4tRL/HMqwyZawIPx6XHc/JaLdwSjbtzHnEJRe7
rPc4c7yIVBD/5xOHGyEIuyXMZudvkNuG9UPGKS1tJ7NH4pJzXOaEBMXqn6SubcCu
5mSNcF982x/6KmX7kxxuUS84cxkDzgft/RCLg0rI3NQfALHvUbbdxYDF6Z/n7yUV
Vt3gulPbkM6e4cR5ZFWPi7Ywzoezq0KKxVvcNahO0fhpAd/aB2iPFP/P7gDJVy1T
SEEb5OgxHYlUjhYQwMbnZfvlClSRmTM9R9grCdpm9kkZKRHBZeVru31YQXMqyvjX
+uPcBVXQLyGSXE9BVwpmdZ3WEMEl5w2RRXvp3lRZkD67+dZnaDDV3bFeZWY/wNPd
YyM02Shj0wnZm+souvC02XMs53zidpTBgzoswCXUIEOBN1wVMVVQ/biOO3ZsQGXl
STHC8Gp9xLg40Qa/ihxRAPlYF88k+jG/cwCzCJ626JlpvGTFHteDak9Ww0SXRFfZ
ALk135iSSCiWpEcxDrt3juawP2Px3y9HELr4JnnPZ+j6ARLZRlyYIm0QtN3V57Cy
/QyIEGW6/16ULWQIoYO6wjOieqkX2MiWDbiclmJeci3xwC8bqqzET46iKBH4Pb+i
njcQ05ZNZdmKzQ4Jn6SMYA75ZlLW2awBf5uEyUq+osgolF5Es9Y6jxhhuz8PoEzx
M3e7lhFRHxtkKfQuPLLw1jLj+TYNuMwt0lolDvRubF9cBvZ2dD6ZSUxOQ3AQAbEk
NFC6MbU31GcUPrUzNL2xxghaenQLqenzUA2gyNpofGZ1FUs5/dehcYzDpgsUXAd6
x9IbW5SCJOd44CTcWWHt9U+ChQhsiZjENrdz/PRGoGAUY/Mr9Wbv/MvV5SjO4i6A
f88QD9p1NE8WOHBH2xEQRK3/9D3r4hb4Ls40Gj+I+O0RrJ4dKisPEMYXDFEE8DZ3
OwLyRPAeGRaJaWO6HXVfs0676CeoHtclXbIHBu5bNMYeMaxnDtJnhi1Pv2Yf692L
38VWGeYhiwcAjgV+yZlTh50Vfoi+iMinB1ZDZMDnAoLf/6L9wsigdRGxzy8MgcAJ
Ix8riNBkQToDS/260VM6jHVaFkiJGmht0VsK+1UKumTXW2Evektuutce2m0jvWW7
K7FQ5FIJJhf+PJhduOXGwuTtjnAWoTDQDRZxvn1r2fV8HAHDF27wKxM/6fdyq3HX
5kbpkN/3A5/FwJ2iVW5TuvIFWBDSZnpS1oLHd7Ps78ud20iiDj582zzaftnZhyHr
mifcUbP5sCh4Vf83styM/eKtHdzE2U+Q7m6OUbcwWJLUEwZWyYLgOZ5YVZzukNmU
Fr3uSDMdDVSfXQTzze+PlXxW5tM/422sg/9akxoK/47Eko8/IZa3p4M16D57qATr
bGVYhtj4/JTiNSwhiEL11O7Mwbzp0IQw9vvi6iJ5ONO/U3Q8RRLqOT8Muf0A/6mb
lbXLIMAuzdGQOT84pBEr6o6my0Ojvk4RJCtoQPQvyeZZMYwVWzvnORyik084B2zz
0hViSXWHX9H2CISLXcn7w5iKqfAf0+jTU7YIdD7GeaAE6U4so5Mop/u2xul/zkvC
zo/hXucKYl0pt15araCBVQtWS0h8+smSK4vU61kPDPpt54iUxeXD6LZOE3ANv/am
yKF0/TewFGlwHdnJ5+OT0+W5IOE/5hEofhKlUJa2hIRbwrPHc8yRgESM+qtg/mnt
iQ9H1hLdbx1fNQ4Yu4Q+dYDuGo6EZ8al5gNemnb3mhQdZWAryU+T1QfxjWPqq3q3
ixb5h7IltM6qlJt06nWJOoJkDjH1b/4m/bYgK+svHjaR7b/bpmIjOiJSrtWuhKwO
6mvv5vMQAnIV3ODBX2pnz8TJXgx6twXWg3r9+kvyCckHEPlt3r38VYoyVP0Iz7MT
deSfVt7pwuDq9HHIc7MHMgBQ+EJB6rbRhofR5/x8/2+6ohoV9AlfphzsMVg893vE
2fi3oB65xU3Q2W2fiXYWpTyyG6l5qU1zedH+Nirl8LsOOmc15uG2phQWaQyn0LZ3
XZYHhKTTmLknqBEs4K2B4IVIHtiBANPbOHTW6GNtcd17CisOWsE3tFyVZ86HHy64
EgV5uF8BpcbNB8fN+v9y3rPAtsSKXkLgN8+WFvOgqi5Qn1+3J5rPqHHSPC5mXgNW
8gMD7Up5Ta3k0FwVwB2ovyPr+S+stPho3LUm155Zn6KLYWxU4GAG0x9i6J8LsHVu
Xik8V6AMXrZgc/oKoiSdhDLZszW6zfFl6hbdHDOjlw99EhU8Bdj/3wredvutVwLy
8t9fASBOpCMRxC+8UgCMYTzr7wz4/gfPHRewhkFc6+Je+hTi9o7fLGEcSRYFPqsY
ZJhJ8+bfsvEG1R5Sf8OZ6F1Yq1h2vfeLqGAIzgvI4ouFla1OiWkafb0uyM+cDvX0
L73NBR/aUIDKSDVoAAgXksLixhQC2fN6VUPs30phP81SsC2sgyrS/oDWchnzFi+S
3m72mBTNT60bB8iEMXORMdw5UmBpeU3Ty2lCXsZm0DJs1Jdz7/lx/sfer+LXR8y1
cIcYiOrXDYcpgxiHjspooqtm2kG3sQZbUeRphWFK6fxF2ScrroG6yZSgokup/fqR
iU5JciIfaJ9q3MwiisoQFaSpGBCE2HFnLtLncuVYKrCKnwFKefZ7FrbarOAHGJyN
HJoxWb4y6K8vnZ+Y7eUuM17S6As2si2jLW6SrygfW3E3MvZZTgRGjXZoQ65daiDV
g9fWAZZ6ExBhzIeQEN1yz8wp+87nHPTLJTUqF3pVyVhg0Gu+q3QQOZNllDp0LOaf
hso4BxJr986gfdN2ZVWcPdgkTQgr7FWfn4t2J3D+KhcfMtiEJWsQx3tq+G18q7qx
xCOnu3TADsYh/LEe5m7Gtdhof5VZAyFuKpWEME5E+jFnhs7qRuwQFPhtsxKt19Yv
Zo/GNCxs6KHqkeHWeHQBtc5ajZX3zOndQOix7V7FIp8Q5fnkvTjMy65/EENCNYBJ
cRxopNkdfY3xKpH++R8ZRFeMeO0UDHzquKJjilsuiU7SQyVSwRcI3G29Lm+SRhIa
asisEWLQv7D7zNs8ZDHF8WozO4GCdgFDycPuLypIUv0n83ccXV0PqC/o6Qxj6CHi
BitYNNZ0UqcU9+enOR0oduks7JBhyGR7OFC92tiR/JTGrvnPItJOSygQ+pTdj+It
g17PuEKlZH/xOLSFK12cu/z1ns4vKm2n5q6HbUwhFG0lnzsLzHYYDeT3FQ5WMsm+
BiepqtOdaMCSVeB+ga0jCOxXzHxs8kTsEIz9gvK0h1JvFDv43LOSxtMhvtLGQV1T
Rk4QrNpdH+cSsVhnEQxj2QRy12L5PDSnNnGIw5BTZhWODM6N8zkZjGiZM7fyQKWe
L4FMEL6ca1CIU2D/BnsbSHO1X5I8ZLd9kDy4xpmZZlv4t58HxnNQ5oF+X/Dmas40
/d8sNzli8qBeVMrMsGvo8qdRtXUpTxTmv1Fv87rQTw6+D2XCaYh1flWWaEul+hOE
betSzAZdIFXUTla3gL2k5DiSWtqbToYmQhGZRgpGzM/EbclQRMw3bgw4QpmZxbpA
NNqqOnNifEwq6C7hAbutrHmeRHAO8Zv/7M10yj1Iw5rXXZWG6iOq/oR+D55T9Jq3
Tn3zvjJtnRxj+LkiStxgGEd69Kctx2R+B25NvZ9zIhZXjaQZZMNpJ8DWQAs36X92
AqzYKHKgvF/9mOAHKY6R32S15EYcbUwpZdfGuoNi8RGOiRQjlxyp/DlwPOw43d0W
2MWXBRx7wluS4qD39xtVyNz8KTSKzZ1VTgY8mG+dGBNVbo8vd80mBHQ4Hm+CF+x+
zIwcMze4eEiTzOIvyd27bQYkVyC54t2RtZEus7IHOpgO0lk4PrDD/NrOFt37x5cJ
WBC6CepmLJ5WmmYUe3yViDJsYsy8f+JCrK8bQijsJvxOCfnc3HyCoMxPCMJKgvbp
nNXkm6ZutTUQuD42HSqvOszvZrQqwe4yw8iNt1s8bzBlzv7Jh3n+lRWbHww7Cj9M
MWcacy45qZ1ijHBtC0ZxAwPAIi9vPzzOLd3p9NjTygA9y5OM9+tCzMyUBjdjuWk4
uP5wdFGWNGsGkeljSgwldPCjOHctYqj8WheTgxBi2CLWVdgUzNFvcFfC+xxHYCl4
IfJhX0sT18oE6xccgiHnnilI/WK8tZ7LVezO2vSYcQ7Iq7/hVR512cT8Yu3ehc7p
K6YGcPHuXGogtS7hM+6V4ARlZKGPpaOrQfwfDm/etxKu/9cdz6ijKE2/7FbYlv2B
qVAxDsNnqmsxZkYcvd7DK1778UIAhZDbh8QEOzGehspk8xy6AavUezDa405EZ8dl
FXy5JPkS15vIHyHT2/F85nqjXSD233SXSpS4Wy/rqQExQqZWXVFDPyg09mDQlmJm
N/Ce2IMavwyJ23sq5RplsXEWVYLt/aZ50xeHGNoHxSvYSJT2Glc19jVpM2FPAB1r
g2hN32LOE2jh7ppLdnOjSmc2uu6TVDPyIVmmWIrsTvoxNslr6Q0hJU4/EDTsclTU
ZdpFjKNLO3bdgTfD/MEkGrIum1K1N+iU6kc1aNvCAJaqZiudIJO28nPT0KsLlACO
R1UQrqMi3PtHr9e/NWnFdHBFCg/d+3kuyTtV9L2jR4VrNiFbmNU8/zrTWDiXteKG
9O3V+Og8y+YWRa0mf2HcMNYenzm+yOu1/c8HdYtgA5uysBMhgMBo/K5UDKe74i+x
lrsuDLsUl5abpkuaFox1PC7QGRn3NElWuT+dPzM7GbkxOMsUNLXuSnOEr4ZmjU+X
7OlbqLITdIMSmiz9GvoAxyGjvhimZ49ARLOfUKMo2pd3Cn66SCKeFRf2E4mlyqfO
SKS3IzbZI5eGONu+fTHuhH90wX2Bv77dpFEuB3H8IWxzWECEiIYnvU7/THvsOueZ
zAhxGe/Mpc3kzB4Rb+pKUIqscEGs/jm2BYMWAMDhKC1hM3xyOrObph5RCFBJhqOy
mHer0Vq76p4sBLry6duCbWFJSsxxPqNuTdiyyprERd9WXK655Pr9+XvDh5X0oCkH
LBPUMtrlrzTIvW0ESYPBqi4HazY2mKoxTUdXgSIfJ2unHQHvtz2QuA2234Jynyn/
vNczNc86eQp3HsNW1TSB6fpvPEu0e/0jspKlWbDfMrgZYtxnLfNdrFFnEsAelrdP
rkcorwogrT115BIqIDHlO6Hki4yvdEwBaZYDZPfiUgF6d+y81TEoePWGunK2VfTW
NCwLJDfkuyQaxtqLaPWtMvu/3XGSivhW3Jtp7fQ43j7qKrCGSANrBEVfVu423H2c
x7fXRhE5IGH+luFD1GB/Zm+J5jYt7qlnUIDaiILKSHXrglJb9XyuI+jIKMwWUwy8
weTkLhMUBfQ3j1Kb6fySzLHRM9MzCsXDPGmXxt1AGt534JLL3R0N4g1noQry+n05
Wv3Z8vPWofuzIHB++y5pQ9kD/w2nTegKvQyJVpM/9s77I5tcUwrb6RYyknrtpC6n
L3tQxW5JiuV31nMgdq10EOBz8roMvbsanldXnCLOg0VJAa0d75Gisyqhn1zKbj99
Hv4iMEJlZdXs9gOQBeuMjvtktz/Cx7BU7fRLaOagVPMzBBp5GGK9GoB+4+0MllvZ
k5sNZH9nFZsHwA2/tPrfHr3owvg8+mx4oIVWDTwlrOhv56Hx65I9L92PnyLLdOpp
0643dTTa3Q4uU2Xd8hfQXMH9J/a5I3/XETMPXBKMEoMbCAnT/5jcPYiPuBb+pdPW
amVr5MohfmO1NSdoJsofXJPl26WLNEeiyQwwu6wSFH/sjPUk2yL2VpyppBUHrmf/
yuD6kAeKHZhwrXDc3jaRBRAHe9wPrV2Fd4O3HTiDfNUf0M0NyLk86ty827LVb0K4
y5ak49uRyRLqHT/5xFIFoiWrOP/1VtIunNyPawiRI7HEDGAqKcreu/Kcc/kOgyUK
bxR4pcmktpyi28/i7pwlXxEhcN0EzdHCKeqlLguF/grE5ITfBGfRuQaUS0ThTLoH
qCvPfzQ6Di3YR8gW8VZ5lwyGrb+z8TKVHsWq6jYnDoxWt7PcPLS5Hu0AaUbblZtB
t8dhoFzt0OSXQI5U4CCmCze/flTABlHt+2xHCK1FK9eMrh950XC4t9mJi5Y3UQox
mxTD+fBQ9f+sVk8qBHAPBNpqSSmRwHy37xjkC4ZwJv+Twd06YfPbE/MN7aOm9cve
JjAbrZnQ1orvLdWZkIvq9HzqgwR5IiUyNzN8+Jip0ruExNpHM4AMtl8SS9pgXcQA
x4GRX2nJerFv0toG5Hm7rvM+IfOsaNnbuQJanT1pemIkxM1AcvcbIJBMu+rGXv4r
e0UcVM2FqshecaKaEKvNbEgmy8jPci6jBhJpotL0wr3HFbhz7WDbm3wB7RhdzCyX
JkKK3D0oYQlfKku0nKn1DZRTKk7eM6pedZVOYya+VqhfGoBMv3lKYXm6jpRQUoTT
uwVdbLvMPY9ct+qvWcZdZHuBdtDFHrkk1cYqcBlKh2OFccRlECJsZgtAsw46NMo9
6GwOgLDkhRRw6EZqNcRxOEeNUh8Kv6m0y0KY9t0cCQDY6JNiquozYfS5btueE01u
F2ZdbPqirzQY2jPo74mZ3Zpwyj/sz4hdGbYpMT1JCV8x061ZyhkrrmgaFe02n0QO
8oMUVWkASpjILoYTubq1IjIEva1a905sC8HdClVkutLzyHV9FjhvA+R5wjAMQ2eV
7/aHBVxnGWXLMA/mkNNZ84sUJiVdKU7YXPdFeoj0rdQk/6APf1AmA2wQnU3CujlR
bjdM/+2vqyDrnKcQd/xMOBiutvzkt2UB1WItAEDOLxiW2nPo46ZQizq31/x1jrhO
m8d4uU+9g9Poqv+P/4eVzjqo4g7Mo58i4dp9FxAlmexWOyiRPgbyWm7Okn6UW2Pz
ruzjvCj21HdTYgvq1mdDaNTTDWDTOhFxXddUeDG9Ze29+r/MNAeb+KwKjhJmFJ7+
JqGdB2/2/iAbTfRoK2DDHDlV5TFbFv4bkRIH4i6k1gKFPf2Cg/wpAMvIX3EOaPrv
eGfRhm9AQg55dWuqkiNT/v+0vqarRL3pgW9FDWKuCp8Gp9iMF5bSwpyb1jm2aqdc
qdiarcp1OIurcORZr1IrJnXaoYY+ZXOKYerm8Cwm1rs9E64q8pWTIng/sw1cX51z
TTpx13gK7Va9IqsRcgEz6huy+fEj8hm1MhXKYZAyfixj8iJ2tSBLGz0rXk+3xunQ
gEJTA5+29TN6dGqZO1/05xE3DY4Mzt8cpfuvhA2ls23rMJQ1Nqf3apqBGKmFupz2
1EuY6iJGXsfkQSzx9JX4vJPbS5yUa30YBC7Jyl0rOWCxv5zoeDoQC7Rnxn5L237w
8y9tnqF5F5RPnUWpFD89SFKRK7OkXHLW1STpa9H4F3McyF1BfH66QKxTbzHAFONR
Sx/W0mCKh3UK2D4R0v/1+cSKrPs14dcgnTyz/9DHUO4dow3xtIwpcR2xj2k/aVP0
UK9q9r99OL4kWGqtJ7TnHa+vqY9GJ7CyEX07dSFf9LNaUksTSYPSbpwo6L06SnVL
R8s8UKf+yL078EwwNXbnELN9AW6LQKw6dUm5ikGxgb7JGav7sqk6mXj6oFE1ktiy
6lqYiVQF07WbJPdgh3OsYTPRwhqGwKYE4rz0j+jthak6ow0jvYvisceyGDJwVIdl
Z6W2c05AxGIcuf2z6twvR1HQM5geRIYFlupxd4Ub0JUGI1MW5UjMLlxITgw2U/g+
yb1X21nez9/VMl1W1S32AyyJw76NzAMwkpcujyoQceHhZai1ZM08HyGpA7x65mkJ
1yXccqjJwMiWuXUat1qcad/Tbwn5ZSIBZ7lLMslr8UXFF6P6VJo61uUsSPuyf/6l
BBZtTkoF5AavhQzpYT5GbqzTT1sRjKFByO+drfgu2I1DrTzg9pSMYNJnBtZXM5O5
QmAcaWPmyenvq4nIBOGDYL8qdZ6u3NFi4fXTHdvPOIv0b+/vZtCEe7iH+kdm86FN
xrZPbwZPngCvmpY8lWySyx3wHQjBIFWcGJt5H1X1zL7Has/sLFCrsYp10ubVl6VJ
eyh5CLMeuO/2dUGexYMLLQKKTrw5BftykqxgUKY5LcgwBGf5VFMhENNorFA/iYhQ
LL8Huga4l9pvrL5iJ9tR7gVme59tVOYYIYSQtvi7+2KGYi898QG70J3gbK4Apz6R
Reyb1EaHffupQ17R62HWZR2ppEkXf7mCdp/gRGx3juC44DMwNndklvMYOWFXgsod
Rfps6/ZsRV1EpSJbZp11RG+ZtGFz6l9cD7ZWMiP2TKL7cJOSZ++ZkNly6FT7FzeM
Hq0ZQWo8Dg2aWt1Ml0l3QtLAC/HFqVAw4UrsWj5tid9HT9YY8j+xkt+mVJBJ+AqR
EVOyaJXLI7iYifPTPe2cxUZdikI2GPEa16ofRtgUyW3DIlCuBzBiBjquzLTQ+nhw
VJYGE8jvb1DItiNfdVQZcQM9dnF2RlvxUJPmAXrCC94Y6N3BEM5dsOPRNxpbFDUr
3dRCgpsbogBmEE5CP3pubdadIw7bLrrt6YusmHr1V1mU0jpgfMHUoLxJg0Z9R0HP
zZP5Fu10zqOpEqTKNz8qXr+qDqcj8AgPJC3nHyZ4+8r84BgDPiHiCzw203NYE/5s
/fyMv86pg4ZqXUN5S21cGiFa/boaHKxn45d/PsVvUIvu/yv5+6X15raQAlZv7UQA
whIBpuoiJVawmqu38ufqGorAjhch4FWMrDzQ5uTEdDpMRWJ1QaRK62FQviv59cxG
V/vpy0XnntsdKFqwTIGKLlhQtbpXbzsDe99xx9mp8tjSzk3EdVmEy0k1bSx24XNz
9VAxiUlSzuMXiNE2rtC9PtSGNVNyDdbhrTPfswruhhTHSwvOJhZCO1iMkA1Cqlyy
fh8n6Hoy0Ka8jRuJgRN8fvfHn/bwtz/xFrH4BRSkZv3WvaHPVYA0N/lGhrRystLl
OTakbKP9xnAlz9hr7M7367jW8Ix3Sf2xIDT26G4AsUMB2tFA8543/yTdkgP/I9BZ
umyMC0gbouJKPZhqdLw8LoxHNHCx3NmQkCuKwnzz5NWyeLfM2leTY7Wn8o2IbD59
buET1S21pHPrlGBW1oB2qc8SP4CHULddc+gC/rWrSOww1Ib9a8HXkeJ0bOgoqL8M
+7KwAK13Mmh+Musi4lZuVygQ/VkV6bSBNiNa6AYhaDHDNzqUVbwhwRAY6wvYXokL
Wf8pBdCH64yAp6O7G9DOsNtOlMQc7NwBBAUE15gyjeIwyVG4dEPvqzemFkYO2NJD
6XGwG4mckWE5t1UWgc0u2Rr/nMX0OAaRaLcbI+lIRlCKR5LXdhuvIY9OtDAf9H39
FHpTYpCcr9R8bIQmiBwUuG47H7GtG1oyKC806ycjknuPEBreXPGXW3TBTzAc29hB
BKbuYZZF+WjhglcztDT/WRe++Xazdpc6+XnEI3CQKE//REYjnJT7jbUjZh1l7zZ9
lVV47W50wDdo6c5mGvcFNTA4i6w+5jqMB5arjDY/K/zfINaqSayNjQDadBrRXmcj
oA+SJSVlR0SYpl1ebeXfJpcxx+wIaLL7Rse9oq/dNsc7F+UgTv7oHKB2VKbdbx5e
8ZZv7EPxVng0ZGwzyJHctDE0Q3EL8t9XN9cA+L8060Waq/98WDzoFRnwMRsJt6nm
R/3j3oGy1WqvRzz1ytnMuhN3Iq69gzMy1gEU0Wt+JQRYZTfY35hVdZZvblbwiuRM
K8NgQwyMNREG23WOmUIIII/wydM0MR9z5EiqykvhjPVlnQsabg3jnPIGUWUGgKlg
30/y916t1Y2hnRdrvSO+l7qjo3WuAxdLpjiC1phsWWKE7JsdBG0ygoyea9zCDY6y
rlkRncckQ9uaYWcCWNw0wJD0Ihs/LHIaPNApJpU+lSXpeafoW8QQO/CWq24inldR
fl5Hqc8pYIsTWZarR5gQT67VuB4+a2yiIyI0jTm6m5C2zZc2Rx7XsSbryhZMkAcg
20P0mt+/M4OxakGlkrEiZMfvZnAAVPUdaAktnY1CjTXhdmI0+16Qm1PTwvn6jbhQ
83yZ9rpuuiMCvo2zfB+b19TgwrfDj+Ll9AvqV/3pK0DNHJuWSrgFfULpaYOdFiJJ
DTqtppLGZGNqXLjJ1wuCLPMeBVOcn+JqOKrD1r0OqO9V6/CrdrrlKu8wR026rvaS
j/rl3LkwaQ3a1KFyUPQqCJeWAnP3keDPeF52mBpzrE4NJkL4Kczu+3l2CegCLAww
IPWkN5OP3ZqkYMm5U2t3qU6gDaC6xB0+hpc52LplXP9COorsW28DMFHphLxZgQjw
0XftCjecAh7FdpiXh0fh6ymSTCPM+yw9nCsM5kvmdAQYxexUWjt2jxMScu/4/fAQ
XEWj13KqOoBn5NUap9ZNE44dQi7PYt3d5AwxpLpLLF6EMMn/eCnIZ8WeeNxZPVcD
j4nkSTed8NeXNFMYRvsuh8yxuZS8LET2BioD6UFrvBNdszA+YeDw2mMt9BMHzkm2
3QtdHYnRnNYARmI/w6smGSVXDYVNADFsF99um5OvCjd35qLzL//O7zUvihmNhU7X
zDr6peVsZwhm4Iw4l3ZWIpxMCCBBuO5X4MojTIsYOioWFL3xvJ9NLsOg/BhY4TGp
K8lK4W8+5IIBExl7Bq9paSgONVfLTO2xM/1eh0NSqtU62RMaPZVNI8ES+MAVs4mg
6YMQNDqmF3nifCJQISZLUuj6zoznJhRZwkl0oViJXFCkY2E3tcN4vkdprASElfJI
ebn4BEAkQlQmITLiT4jdpzvmgM8mI0nXb0xWobvLp4h7mJ/8XL+XUvT3N+v6ZAjY
ICRvpMKs+xrT453EbReIp5AQLhCvXJYMtDqAf9seVHtcBP7v4NC7Bz8Y1CqWIQbe
M32hNkU8IMdwiFqRPm/3aseOlY2vcwCsGBpSvKs62DhehNNKdKkbVQ4/kUoeEqNl
UO8AdrKQ9OMY3/8pOiybE6IopEwsIJjdoZh3KZazr7HSjwWLnKT9CNsPtypFW2x2
6YoNvtr4EOF7DzZkgtVgnZG5t8RpX7az4FO8X7D/9lOANE+jw6kz/UEULUViuXQh
XNV2d8arlz0Q5yOjEF0VP+UwiJGL9fCMojgNg/8KKUqPwIkwtOHvPsZyRzDbejBQ
ELN/rDHBbWl55XsFNIvnMB8x18EVmypzWvltsMnGG03Lz1nU9aee8dTkmM+MAcdf
FsHD6Hl+6pp0XMyLMhtAzMPtyEIcrQ2qfWtDbajdLbmq+18QwRXTdrLvarZUj3n0
+NFW0Y6R6P1Nb+be657ObdelK6yKTwhCcxMPWqBNsxCSLHAt9BllctvJsssqL/Gx
GnfAxufuWCpNFcZduTnJeV+tzufu86a15rJFdVho3Ule7Ak9N5D079bPYhQwHVrN
lHkivVrjBCwH/JD2d0TgaUsB5Lcu+M9TSQA82TDoERm2lDMOoEY4XI0w7ZLbWK99
DLXsIMlMbQeS1QjG32v9g3qpkiofOCAheCKoPSUUbQw9vJRtFwyGMjVPXLKfbJCa
7XvS2QP9Q/w0nkkFR3iDb+L248eQrs46ydQhsqAi99OVyEElnHVuWuF6vBdfpeWb
JddlKocKzNTJl62V2KouFiXuyExRv2ol44ZePWUDqoed3jT5QlDmxyZjVt2TiPSU
aLLmFbkvGVPqx6NyJsahyftfANin7J3AVqFktLjtvOcPPQDuwbRRBXj8nMkoE3j9
JCdK39zcf+jWVHeeWKyi3uXhFcA1NERZVrMzZe0JYXoW6Y5YrxXFGtlHGOJNPkLT
tuhlaLjRZtSPGvE8lQZOPOm8N8HJOf9K3n+PL4w8j7brB4pwUOnxDfKZ66hR9May
lQOQ4chBvB2gDvxldfSZC+W7TLpCEWcfJb6+/iQT1GIxsK1sG7jotPTeRce2oG6Z
hUUiPCWE7dUmxFabkRnawhPr3sYWB38X7bNqxjLu2gXHvJ0Aov2RpwrT0TXPX+0n
b8AWzfvgOZKFP0G8sPvMTeUkwUq2CUFgCmguUs8mgESdexxQLUAQ4woxd2/eRPit
tnhoPa1MJ7PSwyubm8RoQUxxLia7hBIMPCQ+OqL/osMuyFM5Lma/pcRd7XVPxgzA
T6aiMNrKn2UWeQD7J0mIqrNpUh4RJKkSK4AUOPVXVO11MvEjGZXsUZD3n0tVrWfe
ULAvDJoMYw0UTU44JdvaJByQY2olEU3PWu/2p4XLXpCRA4gk/i6GRFp2GOvs5H3U
vj/+tveyRfu/4VT8lO4HeaifoiLSdEYCnoxNTGuS9iC3Hl18hkCeO5JdOfCcVQ9V
e/8uXEb8d7gS3JVX2sEOKLZo6lbdzoJK94gP4yO9TGbqbYjVyMu4UB/nUb6lZR4Y
a5hUdJZiJqHYToMhdvx275ZH5h91VTyTqxqnHpaHCBVScwZajQ/by93w5NXFVUbE
yF/wmYqRZNOSHqfAYAoHx4frKU4W8l6s0A3S0koG5YwE7KMfctj24NgoePRD9/9W
1GrnjPtcR+phIlY0Fl+aLFGlrZYWLKCMxxmIZvQetHg5hxUrge4eOSUujwN+IcIh
NwvQb78n6cLQFI6tlhcq4c9GNCscXQamxtxKBOEDlmLYTZxxwv98F1A09JR1OwsB
OyX6W0F4us7Nk1vrucbEuwElG/QFOE5WwgVrSeD7ohq+lW3Ts5iCYrZkHy4GATMI
wqXwZl8UMPjElng/fN1sBwf8/knwhFiyPz645PXM570entPPWhSLWSAja3PeJR06
uG6gqi4a+1bDROBtw2Jj6bMIYw/jmG5HRxCXuSLZ6RBFFG67DfkZuUvQQFuMmEXH
Y2C5+mG0okLhERlrRC1AmKSnxANp9OVVzMuI+G+UFMeKrhQPXDJLZUUXRYaxezcK
c69koz+OJq2JBAULEYZgR+/r68HHbfIf0oP+EHwYqekWlk+Db1aK1EE/GNdhm1E2
mxxvJ1s66AL2i/mrsqQRG6PfNWHlH0qmc+5WUF8XdDpajyQMB7X9RuRUPxCXV+aN
j9pVEdV+1fxhc3Mz4xh/4VST2zwesNMynUiuSfF4yh4w5sUMtwWZ/L+PM6BsLgJx
09RXSLV3vqBsCnY8jEA0Tpi2B/rEGD5ddGf8L/qwVd8dEQtJOB9d3CLaa/A3DK59
wbRnASbv8lZp6pcdl5JYsQl2VQZlxqocnCHfPR+9Z2pG5GewU8KwVVdKobea8+vh
vCi85oRzrjRIZ/kAQZexYKrgkiE7PYQPO+howOov5Vfgao81g9RCoyCl9EhAz8J1
dRtmc1qBpJWJcVmFgRBfpE6odR0C5EdyVUr+PrmAkDgbcJGzXHTsMt+a4RyZqane
85qMH8ehYGvTRUqfaflDXRO7+Azk5aOrfvPK7XnBbsZnpk0ZPjxTyXM3FWaDNM7h
9uvAEa487ODAD2SqsMvL2zU28FP73sXhh9Ow3bJ3aRcvRrTWEIELllXzCEM/kpqf
qkC3Qj+4UNfZUURxtQVyg8vS83nYroWsCbGfzxkfVG1+bnVWXh4Clnv3tj3khuEx
Ek4HBK61QKLeoLI/ZmylV6jcbL2SypMEb6EkeqzKPDpGckdv2i2RUGr1EbwXLCRs
dZulUKxyYMjRCEScSoCV6h/XWsKXdYThO8xR6GfJaMBsqLgHbRKz6aX4s9Kr/3Os
qaDQt6UdT93NNNy+70EwYyrza8RuQOKQVIheLtOQqHjR2Y7xRSwGI4FivBiMdnUx
8ZkYJljiWX8Ca04owUZgfEyYY86fbP610Y20twxUKT8C/jc6yYBB2YHOTo+Ms+wl
1BJcybAUyGF5I/d3SoDuoLSO6SYrM8a4nM0t/QEoByQ5y+//dRdQWqL4GqbAXMwU
vTFv77h58JnNDPwzV3ci0g0ih0EuEWgrQpHAfoiZCjchwP8yAaOap6M4ggy4BRxr
FMM1Femu3tZ94BzRga+LrR99UGgAxOcLEzCU/vddfBpKNYPmAH7ukO4NPI3P9Wxt
NgZd/Ur65Ep8q8aeXo9PpJry7BIE9laBmAmPwc8B18vbdHZZ0twQF74K5mEgYzdy
uB0NF/M5ly8P+tq7w81yVH/Xs7Gij41m251GzxxMGm+cHc5+n/ILjBHw6nsqNI9v
WO3KvnRR3wumL5pgnW6HCQWlYn2f6GB2T6R2JbGQ5LAXKCDN/AMHwVwRd117lYD3
Qvq3u9z+quJz+3oT9lijN0cIbwKF3bMkAIM6X3cazk3FYvS0Mm7ZADc+/xJURaJC
cLgWpl4Ly8NmRd5ZNNi+82slIfERkU7vV5BiVRV4v15j7KWxGJh2XMLa9n0Omcoa
PrXj2a4ZHRRhnqvHq7FsWlfUDX3Y5zLKQkwNss1jlm60mBLBjhjecy7WpXiZ2A+3
+6nP8hBMf6/MPKMwTXu4e1JJM1SDrj0Egx/BhYXE2vQLsS057lfjLAjMIv8AaGEZ
B6M2MVLVgBU6LDd34Lfo7LWS8eHSgSlaTo2c8jK/3jxXrdBVulSl0bm3xxrwcDO1
URiGnQ7oFm7SwlKNf9dNdOFS3oYNqf+7qrv2NiJ5WTUVD2ZwksQ6XgAUV+G1C5ur
YoI2G9yOnn1o3nHZFwkF9D7BjCqGkMyiEVGJomTq5jkJAdnuZ7cIIEKTIvschzNi
hAqdzQoX7Im0Kcqq8xdn6buzWU7t8hMEq1AwQ1UYf4nCuLUTY3FOS+R3KsQYVxkn
FjOMxZmCQhfH51uQKl8+Qjph7ngXURM07cDmMJcUKK8ojwrsXsfEzd8yHiVWJ/3k
bD4lTNyCudTKfzThmp2T2xXRLyTCWPQGDBfJ/jCAuGrMMylyn9bPlECBuvqxBDke
U4BSdtSIwqe3JPMUXHaxBl6W8RJ4R+M8EuoXciGiKY/FN1dQDv3w2rqptKAcNN0N
`pragma protect end_protected
