// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NFO2ePDigSju2fuz819HWLp9GUDvEZfHOcqHXKi3Ev3Frnca3y9czGIQQZNWp9uz
QtN2hBJv+G6Qzd522yhmSdquNiaZOzITk7O0IvJQy2NAMOTWdRwXwlgtSfLKixMb
0ypaQnw4oG83jyQE/m4Q66cYMgyYQ5scWA5IUVzGzss=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10208)
kVJtIM/mghGEqrWyN83Tq0CzypH0nyvApo8F8oEUzqC+2oliaOBqnjoefj6dzVSE
rCYmRsD7Oz7m05CGeHm9z+lU+ztzuQpJg9BICGYwB1RuWX0MQK8gX3rIXlRVvWVe
NUyvCCJmoyj9o7xD920tPsXPdC+MCAhnT/JAaeO/ZtU9nE8jceTIZKn7/PSn/H3R
3s3sGs3IltHNzqHBL3AX429x4A6duXHJWGdFKkAB9jtttPTRyb6yW+ZBKZdFPT5J
7VhmjPTzbMta8s9zh8ze0YoQm3uGmL7VFPoj/gUzpDfmaALf0N6YFs5ZiKu1I4JI
1Avf2w4qPbzudDhh0CfeQ5sIDGrn9rW+vF2vEUZv7XxTBFVDrRyBYfGPW4AtEwB7
iqpmy7c94ofAgBj6X1SiSV5MY7EEZys1A42ETae+k3DGdJTNPgbceECrSo1R7GXo
GwOk75v2TJ2pbrVV2AZ84RKRZhfQUXPd1Daro3EzWjyQTkBIudn45JB0kGBnuKQi
kFcQU8H+CrbGLCzEK6XSbnZ91UKi5MD1t3oGXWHpciBPlsHK89fli5X5OgLOxhSW
B0wVNiWmZci5/h7jsasIGA1kaYFKZmrwOTbNOyMvnNeX9wvkCeaVMhhIMPaYGnvE
oE2pT9uQuylbGE/MWqcLiNTIXkBb++zq0oRdVV8wcFoBbt0xmCinpaeclclnGqMK
wxD0ca5o52+rsDaV01v42GMBE5+D/CSTRmN45CyJbdO3Bsf93WedOjnx1xNXo4QA
pCKJah/uj7Rvon/zKQpEfTLZI9AVX0Cz6HT+vlpMdGISkdx4xfcW6eG393Km/80v
dOl98nTAWpwfHRGEG+meA0tsNtqsEdV06vQnJM5ileWQViDPU0h6Dz6zZKo87BBS
WDrxAH3ygcOjKbNTHtok2U2Q4p33N28xEjKI4L9a9wo3p62wUAVRFKnfzyal/za0
aAB5IOQKRWmIfos1Fde6Xn4fAT6ITv3dqdlxJY0jd2Osmxfqu9l6lLrhNQMnFOWy
zzImsPWAHqyLN5WKtGnlU0AjQrRIRnR12rqt8IFVdM/I8+RpSJSdMyossJPo7IT7
9LiSO1beh5wji7NQbJcNlEkBzfc6PQ5VFNBflyFsno8clU97hJpvnplHR7NFVHGf
QtXB1C/amikzbHRZSlARiPFBVRv7YqCRCmLd1ZHjYUh7v3HL/lgD3eWVGMl9NOeE
OurYu5wgdFwa/2EAi/4VZS7pwrjETb4piGB+OrqWMT3ibnIdKJT0C88SzpIH9FFh
saRKx/hvzNwgKUKEkiLMpkHy37LTeim6fdzEkjw5EOgR99y4iqjffeKCDe+o/rG9
Qa6HMyge7Hu/WJEUGtKZLHUM7o4QLoLf7wKP42E+tUu46MXcLlLikZYZTKE48JO5
66dJR8YJG9EDUYc0f16onAR6ywjRi654VeF5tx54bd+Gr9YtcUgZHbL0B0mq9Qot
kdLOuxMLhVaKDOBJkjBd394swLiQGLMp3avarGeRpR6qtjPMIOWxQ8I4Q1+OlA59
k+MIxKWZ+/CHKX1aV2mb80XQ8tT+mBh0rUFw2WUbCfQFksJCya78C+m3BAx+a+vu
V5ODnOjfjJwr3OSYLHG2gnj7aMtrn08qkczbooNYQ1Mg0JjV9walZmmlS3lspfsn
wJB2ADw71KzR5VAI04DIWlFoEJ+paMP9cpFHNwmZFyY4rNKk1IaOQr5XAzpYjRpX
hDgxWRnbFEm1IVpuFa9y6Miwg/qLSNKLOP67Ci2uC0vfqj9xqeKElCa2tQNnG72k
HzUvUU0E/0g8vLiEP8PZtgn5PXIz8NK8Q219wRnE7u5ujsur5xsSo2p0a6BjVCJ4
Sb80Bh6gz2mlmUl3VVDtB456STi7d9pCJnzIFa+QX+7b4IcCPbFVJ8pKSCxztBCB
XkNJjrvY/9v1GlE1neZMXnUWnnA6JYQ9KgQtJrSglGN3OU2IZsMLH5T4KCbmaJIz
qHtbolbzx5Ujj060lUSK1LoDX1GYDxWsX+iczXQj50JDf2CSDeW7TNN0fsRKqZ85
kRod6nZEYc/tV5nCxeYVE7nTqIeW5YLav3bNTaTKeZ5igHL9+CbOvFOEhJ+Vca5C
l2q4vHCiJvFm64/tJEtgEzIElUAs3/2NR+bAYnkYuLfE1G1kUvoHVnlb94+eAxkl
AiMZhU51Bq/hjZVV8B/C5rxv1g8xK/CmlDP/mD3l8gvXGWAzeJubFhpnBHvgVDnn
oHuT11XzoJk4eTr600RtpHFwMdCII0pIn5oYM/KRTBZocr8G5LeAQuxzXVFOFgv3
N+NWRNGAI+C3H/U5Gr4T70ysXzEEY8fYBw5l5wICGXClAGDfevUl55OAHmyyAC6x
6d5GwU9pdKodtrdhU0fJFAYOo0XgtUWqZtt1p4PSnWK7z0wwjAyI4XegEc49T9iL
1Z5YjBuaKBEaF/Otg5OoGG94xk5uEDChpCrfObx5f0PUMTAzDzFGuWaR6WX1UmIT
e49j6lEEaBdCxb0jIJHWQR+Z8R7rd7kYFP4TgCGC/UDEBNySAeXIcGxqhxX6etTm
VlMtLJoQliffQ02heUfPMAwFH3ax+p9cv260cy2pEb57aN38w1CKf6OAJiofG1m8
Hs8So5fPnv/t5pCUfvFTH7CmqSPt+5AwYTJXFQnsk8PBhdobxHdyQj8IeAXNBt9/
n+Cjyf2cqkngnWyQlcj5dSipIO8kXp/adl0V1FD5sbn2gN7M2MZVBMVJTgL9XI56
L1xDRveVlpKz6HawwWk2KlulN/bMMoj1uktt3QBdkDCi/8jjawV/JRI3RHJcJaci
4VHBYfIC7NObAt5qaWOxxYPkNBAg+VaUd7TANpTwr2Buuo1DyLs+IEugkIjFGb0v
olpJaGVjsDmZZC3rKygC+ZHBOukIx8m/fIEBhjE5glrHNtAf+ZfFMbzmbmVmKgMv
499fCiXyR7UtBVTUb7VgcGpKLhiTMsUG0bcyTxnsFtU5nAztgZ1NttBvIck0jaSg
FWYAoFNU+5HXsyhgXiB78MT60ZFoMEv24VKboYg702o4A6CShqYf8TNzbCky3VFG
skY8ho0ldCJFZx0GysIgBIg/BRZQUaWABvUNVXXSBp36uvtbbmXmWr3E29hIh+MZ
lycsQBDXV7nEwH+tYgLYXfEIcLR7g8x212bQ5fiue0Cd7RC52TaSzzXbyytW8UMJ
Nblw0SEUMFoNslhBv4TOeEv3RtCC0JPDT7ZX0QIswl7HSVoqMuSBcibc6jdhH5dk
o+NJanbyokRs2sNTFb/WpY7yvfV8qMetqWd5FjUiQPj+1/fYBe6eFWyiM6AMS4+H
yqgBJfzxdrSa3kwdrn2fuqPdoddGoUcJ69DZSLXjyF3UbCdozr7W/5ROJNEtr6CR
GLALeyF97m+c7ImfcihhciHr0+I/0kMAYEnbXWBVooB5WxDplbuBKsIyXbHNY+Uy
5FBbsvemkiojgpXvTmoS/040m7Rb9TID5CTak5FVgwIn4QLLal5X87l4yH4UuIuj
hCYb8xDzT+MXRC/WyPOnDOxAbPO5GSxF1Rn9tfOJQDBMzpm4BY8VSc+g7g7vmtaG
aX1Pq5BMUhovjMDBRNojfnbA1n7WR74m4wIPHnUqZMk5CqeY2YnDi2mNOfrEAvD4
88r5W19RcRL4YSUCPn05VOrw3U8tpbhE5I3MFZ8YT05Q1Rcjz8sAUIa+E4gHBaGI
n3u2fE4yoKYq8nXi8t8g1Jxr3pGiuCBa6SQN12RZugRyqiWskcBUGhxzhfoFP0pP
zCw8AjEvC/thpqMvV36QURK/NgKmq5oFdwIIhhTKQCsJNC2vXIW9lvnGRR5yIMYG
l7xcZkKgCvQ0iXoAvoYnPgAaugw7/JmMYFWOnSwFo7Fn9KN6XxuhPx4hSTmk5w8i
0UCBUUS0g42KshPq0NTx6hsn99cgPdMAL5DZqYUg50y2A0IfeqsCIi8GgYIzWxvk
uDz3h6yi5mPsKGx0Q6j7jZtWVhceH6Rdk4J7AgozTO5sXzucIcj1BQ7Hp4XItWZW
ZHDQGRrxCUVF7gF/719WKPvnvcIN56cB3tbW/3vLjwFgMlB84SNY653ACHY8p3qY
7dS+oJu3yHYf345XPXnW6A3wKNjpbvPfVmfjtJCtMW1jla0YcH8JrHPMhQoG9ipj
Qi9enTymwpYApcf9lmsUBhQUudw+yp5pwiVYnW7w6m1aPTWmfCgl/W3AFIB3zd3I
htGjI3KR0qI+Ubg1avvLCbBQrjROHAfZgGKw+oc9rMesfS/SZL/CG26bYQb42l/9
W10PDmMRLtUvMPyv9hFMApvKxK8W2Im/rW7Kq7++5/KKXDe2jhWXnTHtPtLM7ikk
/t+GVRi2dDajY0OtsLoOi/DS98Pj1a8pL1M3z2fp+wbDeKVA8oz92Uf2KG+wChTJ
suONJWiPe3MqsW16Xk9H0bGg73ZsFCe2AzvzyVpVhYjEy2xo1bFAnn32QYTYdiyu
B3d6tR93s6dGWLr6LKidYD5Ldrr/Rrj6Z6X+4Z33TeaOS5TcyvqukseV4poZxH9q
//cErqH/yOT74VxSIQBoDwa9/GLvt88XPvuctYB+o7OcXUvDkZHIw0she+ZaownD
RK3e/MR/JIRAGPdqqiwcFktA2FXBnHkJ9spxAHB3ZD3jwy4AFNemNMlwWo8l6zUu
qn5hx8mUVGKxDKRA1MH3ijnsFOnjVhjAkAL/n6tXDauCzzAEdOCVjictWjrV9m/A
qU/n5/ACj93GLoI7oQS8tzqzkl0Rxn1mRMT7Ho5e/kJ+a4krwhCL2eiJSvkgSbCV
3UQ25brvPrYD4sQbgz10zYWDYxq0FQBOVmCBp9u5CpiixSMb2ws8kdi3b2QnHo6J
JLDh2e5m3MZOluTmYmuFyFv2sol/tfBtx5G/R0UApZmMBoayGXO+BZAZfHX7Ntsg
iMXU2VCAaJJ6o8SAsEQ+bysZCwB8Z9vbO07u9N8VlQyH0aoutBC2GgRwz4x897jO
YAmcU2FsFKBWLGFGqyZo0oEO9BUpCYO5XY5UzwyrN+plflgEJmYub4ksDHH0sYxd
4cvIKggCyHM4Z7e9EJWE6eoX5jmMUsuXn8wciab1xOH4hhSJ4MaLwEoX+Ks1ws54
fMk1WwQVZ1/lpFQSeD8AiAOkQ9s3XPE6MOJ/W6lVZnvnrM3mpyW7CyXYTKJpq0LR
gBr6UBEUp8Y0SCO5/dpNi7QGKfPzVy1/TbjREoCDZHQ9ciu3NfJWFdHdcNRqCduF
yDK/n2DDXa0mBYzRZughfIKZi12g+/asWjHDOACMLzsEyk2AqSiuBOfhbUeIBVR4
CuFsfrr+hysn2C6DvIXB2d+zzesbPdZ7EktRNGK5D9OEDw2sb1sE5XLi/fLJuw8n
0TK9yn2lvMklSa4bjkty/5N3bup95CM7uxQ6LiItErrnUvmxB4HbRcp8Wit/4TfU
uFn+B9BZiqCYfidqebYnsUYSE48ceJCRiXTvoQ2bIsGqmyRa0elDr3aueAnrDArc
ubMpTWrsr67FsbeDqjg8DxC5c3PfgMdc9lctxLNpcWMFhebsR/KHBWuQFxZMQq/3
OagFTLQOgxXiN3bzIK/D13i0GJcR7GeQXMiuGIl1v3hKTsbkc2QFw1Yi91DDzFXJ
N3N4IHStLI0MglGJcKvATq+eWxh5q1obCUCD7MA7Rg5h6LNl8KRiUF/0CvJwyIbF
Vt5TdB3DJX8zAcLvQch/v97eTA3PdSP3Y/4P4wPkk8RX5r4Ux3DphLETvwL1CXmJ
URW6YXFEW/JsDgvdD3GxG3YWsGTE0o8LG1ifdbS/sT9XJPiLVDvkzY9G5BWqzsKr
bmYPAKTxnOTeYlVXcctK/fSCgnv39bucIcRMnkhG78m53Rva8lYQOKFSfgr6I123
lW66xNdzavq7zpXeITv6QRgxt/jPJrIr9Y0sP5oKr3O1xUso8qrg8DM4MVmht2rF
GuLWbuwGijUoEOpQBEavnXLV+iwxBh2rWofZWTtNDUopFGRQk25gwJetV9Kix7/m
tJkRzEfbukRqPxNTdAPksMj94Etu5BCqOKTRZN2g9Rm/HR7IeW0NXqPC4QR861+R
d6OMXXboVrGww2VI9BphRUOr8f+a/nEJTwU6yLTbxfZ1CwmIPMwIVS8IvSclx55N
JBtA+olrmNmoSSUTm1XI0BtYibD77QKU9DUt1U4KzKYZxxeWjoYrO2oo+gNH31L5
GAPH1e5RUKtgDfwd+ykjOb0KjMTQ54nU9iE0upEZhApHCyi3n5R5Xpq4SBGgZLRo
APcTL1vrAJMM4QkQhAbdh8xeEbe8h3Nt6Cu+xlXxsN93PLoLZH5jcnWb36uPy8TG
W/Q0g69yT9Kl1xKQv0LeSCfx7+BCD18tzf1LgGPG6fvkxFCQ+K/rffVn9maDOzEL
wKxoiKlxamj5S/pjAYDYDn5lDWtnZttlSTmwOoEjlfdh+iVRYsON2rFHg5H0EPpJ
A+okmgQyei+NG5wmYi8dW2iWRSaAskl3I7oqbBxsyZ1wE52fkpYa9FS72BP6zCxb
oQJQl3p9e/FCtUxb9L3C/tivwx/AHa7boTYzOKczYmu/55Qh4Pqb1S8nGEJMXjZc
bssdt1RcOOW9fE0PPXL4/aoP54EO/5k+8VDb0tjURIkXAL9jC6Bl9lEIR6PmP58S
pZPdiTk3BIxlp+Gl9TwjUFe0gEesCSNsPZUXn8L8yv6NJR9Mk/YyEx952EzNVAol
mI8RUURAyQI62MR1W7Cve6aH45EMagiK03L5tyo2kIAsRJBM2Zr958IzBqbzTNyg
xuAsS4xMY4L5jbZ12ZLwgi8LLLFB3NFf7sw9PL1vwNCG/KDu8psfV/xNkxNM+bOJ
dofcm6ce4vvpZ1o12E9fQYuRykNhqgTJ0Y/DDMY3FP2RJyQZktUnyT9bGZRGLWju
N4uCAyLGXme75g4gVYsRFNkECLv3IvNm/K7/zieNVyM2x+aBRgt+Ia4LpZKyewNV
PMGO4LwvMFsltWZljZlv1scgJSxlm6b17W+BFuW0vaFWlZAGK5y7e2ZRaF/pdXJE
VR31jIAsgjBr3dnvrKiX2fPXik0irOrw9xBrPSTzeRLeR1Ge4ft6+oljYAeK2rqi
a6w/Rxncwl55kUze9t3v+FXAj3R7ZqE63W9l9CVrYU7OaY4ra666xQAoLP3XBbiJ
El13P9nOd9UQRzmOPNknb7XXL18P10UxvaiL8vPAp5FFlerqkrw0Q9IIXobl0yjH
nlOtHVqZeOqlNxJFXynkxrDDaaop1HBJ9LxBJ3wfd6U90AXBF1kY0U1yxMrJECog
rWiww7903qpv6lGBfXxWZqth+YBzweJMAV263UDAIM/WKlpI3Jg3mE6o8wEulT2f
PjVJjH8tskHA8gm+luNtrHdfSqQT2oQdWLiwbo4llnYzyvJzrZ/Dtg09JfxJ7U8n
qFMVUteNStv9e+QGeprtxkcdeOa0b7HOwgmsBFJB5HQLXJxkUNXT1XUM7Sr99wJY
QYF8MKyplq/GCTJG9tbjU5w8RbkOiH/7F8+ALt3WtfzzTNHgjTCfBKQXWtpl4sCk
nUY/uo4pfGgdvsNkGdpKhKnLzL51Fb2XX6G0HHUaMnwk/ODNe1WiXs2MIiUtxZJR
nXizgJfhNlmz/B4tWcwEN3GU2KIeHal3X5s3fVesTApoL5nUF9IrqNyElJkH8BqS
aeuF50bOIWY7VPvpnc7BVJQuwh555vsTxTRMHbilL+ZTEcRs2fFPNxfjUGl3aWCk
4Ux3h/HDO1LTubxcuLOmMWoqK0V7CuBJ3Iy+zzQ4qWnG+pgVQ7oXykhte5wAgG7J
TwMA/dK0jox1tROcWg9fIHAGKLgTxM09+00b3BvyG9wBk7Qi2CNCmYERV7hmfW0D
9zIDa06NtP3lofNm8bJ6Aux7fK3daCCIkjqSlQ//yb562eTkgFW+m3usBis7HExg
LwVsnBNFmEnfhI5DXa4v9jd4fntMVq4mSwz+taDdNUgc42GGYELxvRVC5wWRDbOr
Y5iz9Y92hdjQL9uHrYCcpOM4c0pz941m/ygsgo6+axu6mSuikzhN2myYcf8bfc/u
NoRO0WR3gHLLJe58Yu3oKWZEoPdntknBTkLSsrr80r/wf1yE8ybkoRgUhpAWR+UY
o7ZYzcdPTEYHmTt9H+k506Sf66s8q7005rN4smpQmFiFB1SS6vAsOcEyFw6xsWTd
8l9WE0sMHUSDvPQT0h3EB3b4QPkyQH64FEYJybdC2EeqyfsHmoeKZCCtKuU/m+AI
IGL23m4jxkY1LD1FpdVBk3Br0YQPS0IkKsMFZeleGFd9iNaqs8UygVyagDn6snW8
FeoVTwE6fswO2+BvTVsbjxm/VxsRkX0bY/bsOkuGatbMctxxpZ+sZau9nPyE1gV8
bVZ54vQiXu9agfM0cSkfoAQpSoXLHLAiOXUUAY9NNH+Xp5eIGzsdOM2mTw4q6bgv
Dc+240zH49MIUGrI3AAjkxlg6Tdt1v9K2oryGnR+fgHY42S/M8v8HmiWdAoTvRj0
Pal0JuK+0gyB9QZ6YJ6mskh7q6t01bja1sqn+rJKWzsuQsREGcmwM+wPN8lRsDV0
C1PWHQ9AezrPLXemWt29cnj/2fjj/YvTR8Xy7w8bNXk9DAkd3imb3BH5ZgZMDJEz
N0HcH4FRZ1OhPBUvXm1pRXtO3Nl3phOpVUjFG6XdVukJXAAm2XEDxjNLovC8DsjU
g8W3Wj9mYA2tHrGPyAh1+hbfSCrQyeqs4ctVaqC26mJyxlTnBiwDG7XwhCIaAs0h
ksb/z5yV6tfsqg1sfucy0O3HkvTydpO+35c9jV1RYB9RlUDr/zYuiyfDASBXrVeg
GnPtd5Xvxi8h7TfcYCFF0v87KMbWKrXToKVBtxDqF/oJzQgvpKBcvYLcNuVlXZ1R
gAaHu4ZufkdUNQ+tRP4tdsc+QIxh7j5Rb67/VmFv+V1BzPYAEv+ONntT0uyRf05Y
ugoD3Ir8GEL2II4K8k1RuRZUrgBxOekyJXulC2RcCGh3gU+fu+WTmcqSNw6xsHI7
UfejQDPvWhurNjNdvMBc9IyoQWtP7rHl2STZhi8r+gLLsZUlkNPVvxIySK+xuKTy
NeqI0TeeEDsz5Sy30nNx1An96ZRd1O1gONWLVubMcOLn2DIpTd+wLs+bbgAxcr+7
KK1bPZdVn5Dw2+raNe6MJRSVgsWrN2wxg3A57PTysYAmF7Fu90TMzRugtGdJOZfV
J/zLTKmyl04X+Bh69XSNxYp4g4w7vWufjaoh4cmGehotIzpcIiUs4ymdYar706uU
Wot6S11JJlCrjbt2mh86wE+pJMutCrMuDp+oMQsZyiR4hinoP5o2elAuVY0r78K4
uh++7u5Xc1QAGGro05Evt7aE8sXc9ClbqWEhEokfElAaR6HTcb5QY9065cqPFrx7
9jAq0Hb7uvKE24TfbwdKtXnSBUfISYfgQI3/2rsyoAuJRejALNNhhL75Z3/+D516
J6xoo49pxWv3wfcW9iZZp1PKeFFqtZGC1LNm4M2r7Wjyu1VXuSllocSX+RKl66PT
Xyce/WpBCcmvLsLdBZMg0dYU98Td4UtB5/NMvdBqS1FlR2BsInj7+mf3PrzxGyZ3
9Lpk0YcBt5GmjqNl7lSK1X6/FSVGnOt5zg0jmy5HIY1gFu9XlbHfeA/7mkA9UUgl
a8vxcAxKkf288tTnUfPuE8aOaezygT3BAFeDm/N+n23DGi3L0ZCfkIsJo5n8iDQ/
uqjOx1BpvAX/+6vURvtnLb9N2w2JK4Sl2b99uwyG+XLCiZaWfI4fFVsPHCpmBreg
p6p60Kh/HB2prM57MN6kBBBmjFG4vQ52+bnpIyn/gPIuV0OIt72IqdAoERtr+/7O
6D2g70NECI3AZ9dgkRcKn/6jHGZ1LaRyatE7ws1nAIPVVuV3uwmcV868vVf3IxTO
fqVxAfQOO4ntxzYEnTT8wqfW+DTpGjB3sek3WiA3DNRTisehr6S957ZlOZnqGQdw
Ibh7wy81+yCrneOsiDDhxAyJe/Pf8zIdT/9NYurVeQcYmHe8Oa+hLyb3C6Cnc7Pd
tU98bNTXmpV1VVk83YVrKPg8hSajr2/mi3+8gZsVh6XKmumFtoXmizHqcPZjU1Gk
kpZCntkULiGOzyt/tyEm34FtxpsKEDF4tZTOM5F3wJJDxrPGiBwAfXZY/kcNQaAJ
3JxVjf1JVmmvYfHz7+cJyc7A2dJCEH0q5YsDCFThnIZ3ppEj1NJWGFbDGrrNK7mt
ITIxk/BNDfOhAVlr7TY67ami9MHJk3nrCYaYGVN0Vupf79kEh4wMuflf5tIWD/Sf
SQFowQtZGPN4fV5Ki9H2ba+H/yxYdFbJs2qb/79j8erWBDSwHgJ5sU35FXLOZIAL
OKPkBM5cRGcyUL0krbNJHUO8hpddbCmqAa/mTzNZrcnBaaVjBBlf8UR+j+PLmtEr
nDpIL40TrDZBpJ+pN50stKgxZ+ru8e2xGfpVZMVap9RUvgHT9MJ36QlpDJX5KE5U
GEVW59toDoAYwv479cxhdup/9+9biPljefoQlaSbM3h3ozGAcYPd1Kk3ZP7Syki7
dfDvoFG8EgfVEiFrQ1JnielGQ54fRTKYxhqYiD818hoOHTcjJGqozo4mUC45Q51T
9eCa7EeMFuyGtBL4iI7M+IacxWQCEkIKc+XPLzpypl68/At6dUIWar2U90HDhTPr
rdUCaRypP41tprgRoJQjp6VjUBZdMBkbkYFShLPN/DhmGfx+5ZDYhR0wj3puy2w5
Kxh+qmoAals6YdrdaFHIi/j1eTz1xUjBHy0JiAy93tLtMzX3nLlgCsmNyy3lfrNW
xtY4JiXkEl037OhwfgoMdFmbgSsNZtMS/5d6WRrQt/kckADLWW+zJq33xpfu/5H9
LE45Kkz1AOdt9Oed2v30vRppR+XmJU7cGctCIxWrPWu8gZOLPJ8XHUsXA92UpNkx
SzLgLdFa6zAciYe8MjsnXgiUiNoE3dkRvnytogJb0NlxeAn6ltPqSnE0PT+oYPf5
cvBW1lx14bV5PcTLWYG2VNxeQAp0ZrkiFOIJ08pZW1SvxIVOlaYD1V8tpbYU9Ec+
k7xdRpsaOuWyodmm1aMAsn9RUdi41YvATKHzbzeKUfnl9qKeYf9KxEpCPwjdVYB3
PQqUBbAkWuaLduvwWX+BCDEpSFLRL8Oi7bMA99depsqW6qL4TFjSwBdfefIfyam+
L//+1EDF3MrAmi0dvkun2BiYoFfrEQFBi0S09bcI4aqYB/bUfwSXc09MKb8dNABY
ve1iMnVM3agcsgtNrp8PKg4SyMFaaStKSaFFmlqtfs/jij3mhWyK4D/vS35x0m33
bR97RSIl6pRa+WrLCtn9LHjx3ej3uEtV+EHfqPaDHy0PfEv0u+Fp0UzNs5/uQ1rc
p8lkT1t4F7cbcrArzD7UCIT8OP2GzTUL1xWOgn1wpLAe5r5oqXy/j7aS0BhL5Iow
tfAQ6qkdVQNd04/VJR2oKNL7vMyTX7H3VQaPmISCCtTIvv3G6iDdnvQ5mHboR8rH
cSt9M0vM5+qCOV4ar82IuOOKQazMsy2stLSBrW0e+yWapxQJlhEqqkbTjfvhxct8
FM10hbG7T4S5JpaB4CH0uIkA/8DiPcJigLczwapnEb0Kcl/BneJclniESaqG8uJh
rK7JDkkITtcrfxZn9SMFE+l+e2f6Z1FCnSUsbvYBWg6Ao8HCNMVt3YGxyRU6X+wF
XZBOsHscPNUZLtz9kDhofQ+/rE8D+DmLQefiWPo09ZwTK+BKiNalb/tCVPadlhU4
xdobKQZFkWf+QO8TKWE8mEXfJYOkAVv/qe/Xa/j70J8w9lmXqOWwILLvcz24vknI
OfwvZH8Z31CQZbOsJhjxyHkpSG4CVkVO5fCggBjIs0DRT5bkhrNiNyPi4+QpjizX
u3Yl5zBQmSBrr5yc5USrQpPTwTq8NCC17NcilwVuSybHv9lmMRBsRbUYi5nk0TH1
VOK8Tj0eoEyvHabHkT09LEcYvVSZ2qTTe0vVaA/PAO/nUXHmosE71Badd9tc3thM
rlnyxKxELXrTt62DZl76gR0d4Yvbce/I2KS3tpwZXlHZcO6pJucCm4ALOVvJHx0R
nBh20wVsm1IgPnrubIFfIZ6UVsCfB8bIwmr2LnCD7x6oGX/9j5UtYaFW4nn6I9R1
t/gWJvcXcJPzChK4uh0qvuAEIDi87BoFf8nPYQRSdg4Uy91mXSok2s/7UqLxyBTM
j/p5wTbbs9rdjhVbHjVD2IYy7NaljWA9T0xbEvE0Oa+XOLyHC9O+M5sgDmrsyYdl
8k2R0Q7CdwE/efnIei+DEW89ns08cTvmuHpK1Tg0UnCzSYrLJkujTPtwwzHY9HAO
IP+k2+BnxGdql7jMcWaa9+6qv81B6Kg2LmhyMJYnP1tO7XT685VX9w0RZI1MGNyu
nSrYY/iQlVSeUiONq1yLTXocSlHBPWFlYmRG7BMbQIkOADedRIQalXky2UsqCNke
4uUOlcac0hkY7plr3bcFXsjwtvB12c8PXsIJZmkKc5Z8jTCP+Mc3AN2JIWJWdULq
pfOCBHwJqYQ5WIhEIvvDdwju7WEAxPVoLRUx4PEk9+14j+zZ7nnsfdj3LSGWtrvH
Px3l6zhH1F48EqEuwI2kDW5zave68pvbx+GYlYw1FKNFuW5jdGeFBiD4wzeECh2B
LvQE0GB8Ul3oiJNVmo6z/ZbvpB95x2nG5YnNGoxsJ72Hr7kYWBdRalsxRPSknMtk
WWBW6U1YHDMHoNyiIgasi70cf5f82+nRT90rKEpdrwN+BDgOxz2mqw+MgWVeXuME
AcbRTODRCFb4o7rglWgBX9bwonB3DdhYBL7pOyNISAaT5ZQj2K3zm/GLlBO0ixPI
2tnsEvxWgTPXYGNjg2cDi7eCzsEkeyMVBbLKlfy2dL5w5ghkYDRE9wI0eVgTyZQO
72zlrOctpC4n+dxUUlAgBLGGa84W7wsJ6V7WuCDXobO9fICt5a+0fftIiOHBVcxr
RpXza1IKOeUorOU6BSRx/lqagYV/YcwN98tfH4RoMcLxGm7wzSraH7CI3Pxnce5e
NjG6oQAkCvur6El0o8GjlsFE+cOzezhwAETSvvL3YCLEvnFabR6andhMq8Y4ECkC
xRpGzbnCB2JFxcML7+bOPOxRXqPIGQmkq/raFTBpkFB/L2CemL+vi4lm++MEYKkM
oZladMMiw434cnCtkBVYwxDMKX0EEzyiwoOGl2SAguGzAIcIC+wsw9TmV1yVUn/h
GOI6UulovvtX7WsO8HYYQpGM4D7psqXeO1ucvtbh4d1VBONiVRdtuPacGjx1ospY
oe/Cl4kdPE4ahj+qbpXxQMbZHhOJulAEm0VoOxUw5O+ce7KW7aOxyr/PebhFMZR0
V7fzw+qgdyK3bPkP5AdLg9CBTEX9mvY7DihLxd1koM0kcah1Gmbp2jBjoM5vuVuU
R1vZOeLixCc/2jQY0vjnPJalO0qyzTteKnpra54KDfXkJ/wIgvllkGBBN0GqmT0+
DQdU4yjIz2U02lI1XDGucNm8pcBbnyMGTUUsbSjXppMjHxbi8NVagFJOM6w+g1kk
d16MEUlnqSWxa8PGuQsEGY8SG+8WXW53mPY2Le9QwdQ=
`pragma protect end_protected
