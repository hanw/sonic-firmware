// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TJk1NlaKFYszUrfB33wHghgHSB+d/M0vOjDn8UJMo/dTdmwTMiS/CAD94tTj8I9g
F9MtYY1HptT4l2ib54/AyjUiWdbAJRjA1/uSSEAVYKqIRUftDzw2xkhQOSReQlA8
/Z6Va8ttiO1u1BtNPm0wUkRI0+9TUBsMXRLsVfDcx0o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
ycmBcv2ewmWemNIdC9zqn4siQGQRBcOHT8ElxsZlNfAYodPoxW6XS7Kte69dRpub
8kxwwZcgAeSOIN4P299jDFxjeHBI/fEg4Z5hD6He15wTmx7NlydoIwPO3qj0H8ws
1wW02zj/McZ62W4EUa9CACZyBBRbWlVtW42ZEa+0l7SudV7RJ5HMgXXi0O0YcRu4
oYxWOTaB0/SP2iaPTYiNhyLdG3cv+zBEkpS8zJQjtQhbvPiSi4xh9tm0md8IQ6m2
ptoTt5IsqCQHpzUWjxbs229vtGwYpaeqcfULo6Xez+92HWiMS1iO537HrgMBw5wC
YS4k4Dn2DU4+5kCTV82ycU+SS9F6xKNLYoGyYUgi0SBqlfA/34qVReKfzLYQP9/h
tdOssR17+h0jJ7ZpLemdJFG+rcIYdGUFScAIA4dSkLrv6qH/3oPR3OzcCwfC4LdN
PS78S6zYwDlJxqr2S5OxRYMt9QFZ865IjKReL00lnFmcO+18cAmtbdjf1DCDJ9Mi
uFwywO7nBeciSSIaEOudJsDdfEMUpew5eEPq2aarIECKbaxYfJDUxbyqQkxPniAd
HIxRB3EYa79zs6L+HmcI1f1AzK67VA5Fn4UKtRGv11OcT1F9ERFps7tcPzTxBfJZ
g4A3rKP10iZovEcXU4MTtpnweuAcY+A7I5IznbdEY2bCdN0ckZ3MTQ+RB9lOpXL2
Hgz16vwHwomiHSLnyO6FTOtbHLZtSl+tphi3969BtWh8+lk5s6E46v0ejTL/vs0j
qTQa3N88i2R9k1ox7FW0jOmXblz4aVs1EvfgmjxUhOZv969BkOSDBB52vhuX2KMe
dx/PAYKsQVM5uHbvdtbdJViQZ70iQpNk9qvoy/5rsQo/3JW0Sq6ZQ46CRESoK0Yb
ytgABCPzhk0eALUcn0PGCBZhJGY2WtlvO5FrWLGVANjkUl0Vi4f2wvI4qN/HiVI2
r7YaN48suZF31CBtkti+nembXgoz8rVNf5erLg7bvOKeazSL3cC1oTk0hIGL0BZ2
8P9I9AyM/X3EbBVGix0P33mHGifKEatuQzzKp3AUdYnKSfZLLZzuXYCJX9uGBwoF
pCrFm1s/tr0XlyBRigyk8VGluIlpqNQISjnv38OzFxsIcHcqzDaKUtq7w/WweTTz
EiGgtvSO5+CYHWZWTxs5mLDvqvyL2havHyln+0j/uL/it5O+syvCUzEjxli0suv2
AZ3Mwl2VQo68/1daK7HiHuyiIoUOza4r3DpFaqqCO6fPqiLsskAB3MI8kepiLIl7
i3G2yXwfuxWLIcAAcy7kA6nCQzNNL0b7fu6uQ/7Jt6ywkKKvU4YMl4dSro0G2OXk
uaRTG8OzApQvPcG9JyOL5dzqhj6qHLcufFPaoMuBMd7xJd/UX6RDkEaVAWIqoK7s
npdwAIUPhonKl2cNPt9rJlDT7azk/R/hI3BrU1YPel2pa4gMSoHwKRqmrFURWddB
NU+Iwv0g0p0kYefNc5T4jd/OeXYXON0GdAGDlZiD7+eoIp1mTKo3X0LJfkgZEEIT
WGtTn/IUK2S/uu3Xpu4F4TRJQZ9xSIo7ikmplNGeGOiO8Eea1yjFGudz0rIdxU34
6ox2xqnS/kbY82OVdhSqWxE9dXOMyWgOtRTLyiPFyUivkyoCDRiqYhNfuE+diJZh
ukTHoECBHuD9qltOPCDMxq409ydca3GmX6ctbmY7i/kzdWQaMj27XhskYzXkVOR2
Xm2hMeXTsg/E+nD6yR91uFd2ubiRwojqOAd7uiEVuE2JeFeUSXbi/qXvdZsuEZbA
TfrGf6BrUz30+fVgZhp4krtx6MiogJgczEI+fdrk4gnOpePxvunJr29MDGRX51mx
oncgUSA5pATQw8U5Ixz0kKFSg6Y+mwIMrmtemBPDSzKdLsBJHHzKxCNnszZbKSpN
1xNqHcwExkqY7jYZjm9P4TMxWvXQuzpDri2ONEnKvTt1HUGiuXGvhlKsCye8VeAh
+UbM9OCTuGLNGjDbaInwxvO3Sx5nRacn9rnX6XCyppWM2EooGaAb+bRSHcis+66a
O2qA66Xwbd7IrMKAuygnt0qQ89El1v4HEZod76mSvRpYlQ4i7v+hEYP91mjDDfPg
EL5/Kw9xI2q1QYdz0NSSxZkFTuYO3Y/yBkgLErz77wxmWlU5VSdkDoffUPvV7Re3
WySqeklevrlZa1DXxFc0GiNP5qcM3FWGbAmSGREqhMUvsMYCHTdjWBnBAZJ0Jtcc
7zeAp1zjCQvMmJOyPnzPsjobJmtCBQMxrQC8tpA3hITNRsf2g+D2riUSTCSoo9Jm
LXMl482e46cRC91iib9d4LcrLm3giwunVLkMhIQkdmxhsdra41uhDcTxSRLqDKzJ
RLSkZNJeyon3yxbn043Ynn8+9A1Zm1qIBp2IQ9jTWwhLNnUjGTIw0SXi2NJ2+rWR
r/VL6PtthTFx4wE0pJRo80b7ud83zia9wSx6/jzL7hVFxWjUV6tnFd6fSpmJlmFh
ui+JTpt1bCzf53r+v5Vftt3HahQJYw6Q0nnbiqkerSABfVgtBSF3XgPgbaytkaiK
PpxyyIUNCKqLVp0UG4P1V26q9uAbzlnEjE7lTA8DWQzRD4uYvR6ISrhlv8NuZZI3
6c5Da8SoGbD9Xu3Dcf1Wdur9CJ/4HGrPnmAZhdwTcrhZgZqi+nglGyWvZJH6gCuJ
E6y3Ck9fvDL9EIgdyqhyT0HQZrkCcY+ZTGLjt+dCbHFqAKakqb/IUV4ig82M/GfY
qhjNmouXwzDvvOnGiTNQFJUB1Jq1c2R7Zs3iO6x6dcYgO9a1dPdDDpB/eEn9Z/e1
N/FHc98WjOIjq7dOD+tQoUt9XkX87sgBqHoBpVCdVTd1zKQpcs8RABefrroVx1HW
4jWRrk+smgVmX07d8C1vd0gouXfUZNUFcTs+VXRDLaP8sZCGaEG4oEeJ9cMVsQtF
yAbz8C7Yii8lNMV2HwQdlzdsyHCZG0A0I23zOchSfSCOuo7352xcJelg9JWe4+IS
LfAjamXTrRUzZE9T2liSh4xSEfsB7g1xixU24ektHkrhCNxNB+piYVfNBLmDbpPb
OhMYhMqhmpYcy9t+9Js3qmil5HHUa5oaXhC6KOpN82xHFYviy/6uZco8bARVFXJJ
SU+ch9RuRNsA5iSQWJUlLANIsKZRW2dVD8C0mYo96l1kI9nJQ0bKG34dfv3b+jM9
E4f+UlI5CrdMJDcZzuXnL7M5L/+c8T5vJGwFkF4oS46KSuwsN82P5JDPUslB7A+g
OHxmRFyG+yxnhq1yH61CcFj5eEajZaNX96sWHVD7FTbHZNpCdSc7/dwj0JV53odc
XDNzUuWjhyfdjUsEMSihi4RfkgGqFRttQ83fGA579z7VI4xSXlwRSW4JY7+C0RT0
skIocxlYwgCSmZkWOkPQiNz3EX5ypXo92sKbyUjJAYxVk5xfmm547khWQQArWhka
dmS0w2xx61TPcUD55VTvx2jB02RZJW+E9K9BDTF5Jzxo3WBS5h5VNb+jHrs3vsBH
DzivTJuS7+2WmT9JoJJghlSxEKUHIDwY+FBCAhoqQOUbQ1zmVS/HFEsHCQMYWelO
XAMfHL3zaNktkuuNvksARhnt71K9GLisc73fk9p8TPh9WN/2llP8SpG0F43XnScC
xZO87EdxKtonELnuIOnvDYbrx06+BI2mavJwShe8y0/Yr7FhCGQOl5wiQAbGeIFJ
5LCeDgegChMgBuQzwMZgnh5cFOTqMA5I3gJWFSbkM7+03J/xA0ujQgQD0bkxlgMU
eflcffYZ9j/BINnzscqgdTKhrC2iFGQmYnu7eVtFNJm9v3aQ4QD4HADD3i5fAyST
3uN7YJcAFPaHkyv05FZQFXLYXlVbqpLLzsd0oZdYfQxLNUsP75APjnkHefo1inmD
Q+d0eb6zViFwECWi/n581yQHV2EtY49GUT+GbQW6SoCezy8FJztt8eU6CecnSzzw
gHNofSV3qmXx/7jPSBdzN7I9GNtzBpWOM+AZB+qCmu/gwntbqHWZnrck3cUFk0eJ
lXLeo7lK7w5HTl0JfuJ0rM/cQ/9Bh471o4EK7DQY3WE=
`pragma protect end_protected
