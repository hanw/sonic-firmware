// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rAHi7URUXWS4ZbqDlvyf8nPGs4HfdsG19VnpWOUbDXAjbg2vTOlnYC4B9iwc2ZR2
In0JK8L8u+7wobSVNOZ7EHghmQ5eaOXDbc7HIOcrycda7bbrKeARPbxrJxmnw3t7
/u7N6oFLfBhQd1cNhfMLGiApPSToLkbgGAvu5FIyc70=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5488)
pzFhPNYJ+gwIiKAS1BjXqXdnEnOw0NK/WZkhJZT8f5vpaxGk0M5RMBQU41d6LdJ1
8F/W18H4QkDuA1zxZnRmbXBCs+bzA0mCs4OUIq7RXYJWe+WdAYP0GjnfjFFsEW/u
gBSXs5ozQpY7plx0zWqR1+vpdRwMb67aFjYWWWxj2VU4i3++nlrR86X+A6ebsBwr
jL3NFwLGw1QbVpgGexaymD4Sxp2s3DrPJ9pxjecskKmnMWoRWq+3Qnl6tLYcXKG5
jcTJ/0F8l/Nq6k1cGi1m9pAxXCVDahfqCS757Lvfw7GkzdNji2u7eL3bwzRQMxbE
a9dHMAtGUzruAeRWCnKMdkY7k+M2HTkPscAvdURZVAnfwqORJlHbGHpFFqrepVU2
5LBSt3Ngm1mPuI3xVfvbgdTnk6wcVgXU+gmUFaNF/eqWH3/sOkT1XKhhDBC6y0Sw
5HXn0RPZaUbTebr2lcfjnw7pgGlWQ0CmiRhpb/duI0LUKxjTpysZe77v9pkCgvRa
nb+plZYgFzIFx0awQuK9pBFuaiYD23tUxAL9vR8K8RevJBAOtWS0SvDiK8irqc3J
zCfhdpwwqMMMp9eA4YwAQ2JK6cHhWUM+mFbN2duXziaEmzJVDN6Dfx/rd2j5char
m9d8ypqRIVQ7tJ7Xyr3eDmbkIf2BiRGO4HiONzoaVcrc8X69KMppQIubMh0gAamI
pMLTeHhmQs8fEOqRONcFuYjC/crP0yqOcdQK7XCOXtslbICO7jOakZdx0Yw1uDLZ
uh5CvsDr5TVjPjLJpvgQfbJAXgmnfOK6fpHhaaVXrU7iL8V03xQzHmppeeZ3X5y0
Rm3t0F3y83Cuz4ciNJS3GFqIHVpnn9BE07l53wL3Slw7RHydioZtbkkZwMHOgJEs
oAlEtE+lN7f8BfMm+are4v7EFHOoAP5Bw+eAh0KsOxNCojkgK2xMh+M5qUyc1kt3
+fbv+Mf6GS6zi/xSQ63aZAHRefi2wE7r8GMlaVcFoaee1636UUJIS+qXSh9egzd/
g+TZu+sfLfhGIX/G80SdwzSOtJg84YtvBXeaYKbiOmFItxQpGxtvb5mXlYdcMPDZ
rqmvW4d6zmwOYeX7ZZbweiCwaaszGcR7gez+NidfXWNDZLqy9QHlDLenSxjN0uiZ
Xix9RoId6ELN7/Zeqo5v02UFpTknSwcbGM1x8VherRFZneP74DeJ+q0JoMb2KeuA
IZebu3zVL1JSir2vYx/kJMaVZfVEBC8NVOwtaKXIh0a3aK5Nxteq4EDH9AzuBQm/
lJe2w6PHoFVDjMMRtEeTulHaywQF63mFj/CltqDpnLPuWSLB+MWD1tDcTQss3j6Z
TLJxt5HYlvZaYkT2snQDfe9Hl33PS7278JhyG2b098KGaB66f3rY6MUxArMgOH78
ymJd1kI6+Dl7EEkWrNMif0h2VYTSOnklqTV0vo/FXRDdqZ1mxNSyNto6FM89MqjO
oqkvKWcpGbnvT5RhRXNYF03TAbu57FloE3rgn+NF6Sjdu+l6Jq/+8syL8bbvkshr
ihUBb1kpInHwnyoCSDZHE6VFdhVUf90Opf6NB4BL1FDuODNxpsZH1rkUyQyQo+uh
atHN7D8ht8PwlYH2RtRwpd+8awHunXorkRXcOVxTGxtZNacuNwlsuDhRjggItkZO
ic/oJ1XAlkYXHepV90nOZyq9KEMvZGX3jdFlewPDyuof01EWp78cwZgMpl7NGyb/
UaDzHBPIrrkTH8I7GU4jGnjcClXH/UNzHtwBBx2OY8HlJFnoiGq+9rL+qKXa29ob
Kym3PS3EJ3zESZFVteLcIZ8n4wq3pzPRi0rG3+lKzdXmaU8Wakg0A45FlSKINYew
Y2YQkKu4JS5rAy+W8hddInE51QESRUVIx2y/GUyOqSD2x3EKySobiezorzzJGtcS
gVOR3yjhjmkWZTBymQlQnH22ylz/5uuN6auimEjs6OYqMT2qhLgkbtnrtyUS8wOj
4FAc+kLKV6ptkkDfGZmJVuKcEXfxgBAm8y0/XbXiAHBWSJlTZX3Xao9tJUzb5DP1
/OiOKT0+zlHPo/dboVUqhQ1alO496TuCv6Xln7NR5YRRjl1KEREfkhpKIfjivFkQ
RY5IDrpkBeBJVW1sxo3GEqRm44K4UezyAiqy47mWtfqRUskrt2wSk2ZJ/qS/9P6H
FIiloXdKMBBrxdmm3vAJQOo+qAhzj16R0Kn4pW34dLBPCGp6qBYXp8LwK4cDGANS
LhnqCq2/3vCB0H4i5FGFZ1OGBWDgygTYO6IGtgKSXVFNMm60eyf4kibk3cWsvlPH
7OdUziNYqTLMk0FpsF9zIyvMI9VBPsKaxfVFjOScT3u+ix8urcewOvRjJJEprM34
Erc8u3G1mRC8tWh8aGhZWXEiM2YKP2jwV+24WYzSoQ/R6xJrEIEHIINni8NS+Qgy
unRMAb0l+quMIKAlYaXxnfQnZCznd+9vBCMGgW39c/nHv6iqjLuKIeIsQarMHpjV
tMCtqoufsfG8NkmV30ITfffl9bG0x2iz6+cRiL/qMitZeYs7QiDCDj+t23BbTJNr
4Z1dld5VS2sCsTHqzgAeD2mqVarlKNLYwEZ7zfGBluvoiQOKfuAeHcXOyKIzrEug
fQkClzEi7beg/hCqd18HLblSkvAQ95fcaJxJr+sevz2pzgm34xdvCTTotmC70iDz
wxlGMMmpJ3G5M1H/NnBCk+Nkx0U3TtABYic3zLq8hsx6qpSRGzk05W4kKteRsfXC
yUD16lUvyQs67g1H/IAqDMIlHpHAjfnnZbXmeQTNxkDujn7drLriF+HwvfG5mwYT
QoFYSU0ZNacfq6hVKzgtAlN+L9iXpteElAHGtHqBBU5vfo5WP97vRmPV7tX8ER5f
C6cbFUsf66BteVLWzJgL64u+sRvNTeN7Gdn+B9N3Xr1zJrs/ZUNd1Rwfw4GPzrrm
OCKwheipP6IjSb2teoKEvaiFsdNUwaGRbhzMzRaCh5nRqNAfZqvYGY3+FDncbgS5
L382i+qQbQ3vOiqbhc1wM21gbU3mp+GE857khFsIaTIM++ba1O54pMT0NYNU37Z6
jKpSPplb5sl0frQUo6K6ArvQX2/L9Hf4p30nZYs/sqaV5Ju+tc9uF2z3RZoFNV81
ejrBmh5vshVY+PxMEQfy6dSDHV9NWV3NzzWohA3ZysNk0y2+OEKXLyer3uCjunUi
afrViMkMGG+jQrSN9sGyrljGkkuLV9OghNiAtY/pe+EUdg4ulz5GlKD315C0RRn9
lobDeRfr7XGW0iFN7YMSBa9pWIwptthXrGuJm+OcWLYdch0kHtXR4grZIdotuBK9
iElaXFCfsAnR2fMu7JAbj0RNd5s59Ygil4cWB34PL6Ep4sMiAFAUWYkc5fvaLiBF
remERXVBDxcHn3HyP2B2MFWzUWQBlV+NWgGVDHJ1v8wjpA5qIMIqXVveV7VCwzJ1
icJHma1nyNel7yvmAmTVdgyfHDBJVw8yBUQHLFfZvaC+YKsO1jMvKzHTuiVSZ8ZE
+CMGBpjuA8wjVAL6PgCEC/ahJBIkWXQ8rptWg5VMf5zbKvXcKaND4reDQ5Lc278F
pqZRYBdr+E8/peCRH2yUkln5BPdlM4X4ddG18qlh3euWhvEIUjOeObweboN6bc35
nbw56HRiK4sqff8/R9g7MwT3gkF+vmZ3vLLB9zLMbHeq8pe/GAxaM+amEM/j4ASv
GBoToa7j2isDWirnbwwgoIoxg1oauzT7Kmz0Xw9TvTxLHeBYm+IA4a4p3xH1zJi5
Go3bZnHPYV9ddNIo32CNQuPBSmdFN8gQoekLfXfe29DXXMr2B9CkJXUqDJ0ENkAc
DiTBBs9+m+pTr7uDbs/vX24IxHBr5rYenxwkyXu7KM9j//WWUPzhh3wzwCvh5gak
Tl1vqcIt5L5wXB/jPJGjrH8n6xLTVJ8pJu1XHy7uh8va7hrvfdmSiWZ9bXx943xi
lz/SFvIWR2AeVSdetVs5zs+hHW8eyK4Rh1eRTD01pm2EkDivUDFql2GdQmIIMdJJ
TcSez2VEfB17nzDwDgRrZOQrBlq/2O1C6cbWPL57Ur0DuBibLAuNffHV9CKiuPgT
86o/yQ4EKWf2vo5wni2pzI7Gi7lzFrXoFFVX4005GuaLOkFlw8iFLOJqtBHRE36+
bJAvOQid9A4XlOQpJ28lgtswyDeYuVNsNxl3tZKM8TYJz3NUmQ+pedfugwmez5nE
fgAeYGR4pqaLZ1rhh1d5sb9LrRcbWvyg81rH+afMvbB+SpjtbJjZ5xC8mE1G9jku
jTXkWSdzGj7XXa076J0kvQ0z3qr0qok/I4qHwUwmAwfgfBg+JBu6pg011x2Mcf2V
wIuxL/cDC4KSx8cZeDlDhK/4Z7bFbvOOz9q0Va0DtShD8b6XqqEmCEwfeI3sRTjV
qqiGO/xMEokiREmMPyMCYNEv8n1Jo/BhryjFhL2H2lKqg6NsUojT9t/TjpFlKTsG
XyTAc8m9wnHanRVD5sTRb/AP6ZqfXlZr/PsuIGMg+/XqEEB+hl+emobDm2snlUjI
J8ZCRPiY8nzLBzMfSG1j2F2xN8ii/6huZ4Nep6BpyiZlRBA5RJqsQgb/d30RVZXT
seu8RLyJDQQQVKufEubcSAWiZNP/iYqx/RJ+gff5jom3KSPOdqoqRktSqRxFur1b
+5LFJM1kCHLmiuvWKT9HZwG7O7P2M2Y48bdPL4eb624qjeqs41uuBbc4kw6OTH1c
T0oVFqowIxsj0wpUv8JlOF8wDFa1vWJDqBfx5UM344HSaySnpuCc2oQI/oe7OaW9
PnzGvugpOq+Fc6aQfOECR34C6Se3o5nYJBz4qAB9RguEZDBnRboQI6dZD8RiPlwC
hKXPqN9s+twBRTAVUOs9m+DKE3OkZu+FEfBKgT4YjpUOxrpW0ceq9FYvvmkXjaUs
d2vKxB1ZFdcbmm2C54CnInJ/dtWXwTEw8qZrNfeY0Z//k0IdXgbDh4l5ReKGYGK0
ZPbZtH0ZYLvLDZ4r5UU61jQJ1/L2jxHbibyme38eRcpsjvtDSJGlAvudDzeNVWxw
qwckcoBV10WD7s0MUn1UMbG5vXQNaZKbh0I9w/hff0M/bKoTKXiPl35pjHR8nrcl
ryz9XU4XfLkKoJsZVj1+N6y4bLXeQ+aXV6gu4zBYzlMcNK8qqaDQzbnN3M/Sa04G
RtxKfck4zK8Jlb3NsvkMxyFdXkm1j/KGoziDhhCRle17mqQ7xb8NPK/sYtD/Zmia
VEjU55SrJfQost1UuQzH5+68boK5rEfCuXpz2Cr6RxxBV9pMugcbU/cKrLcxB1az
CovCkQptywHDHeGeMhirVT+SW/LYZ45a/b5+vQ0TfDJayJnzR2DUCPYmpxNuFk8F
DsvvkfzPThdwOmZqUw74mS9PcFcvQl4H53m5IchowURT4Y9OOcyvpEJRICoc368j
f3hnu0lmEYLlNrHygLuPkS4zLrZE7/XcGgD+i6zE03rcAkBVNZ+GCpTeACKXbVuB
1AWTOyJu+98kI6OfwRiw3xe4n7o1XHY5Q9CzK+8nnRJ/hfNWsggqXRHoyev1udTU
aAsREBSsEhlqJYvhYL6Gb1QT7Cq6T/Y03GsX39Pzu5sxM7+P8itWk4cIVBdNU3sG
4c9XBJZ0c8yr48KUUe9Mas+Tr23rpUI6lbTKDHUUNxhONwtP4ztlFHFUJcL7SngT
Zgkuq0Oxz6Pp7hTphp6/tV2nN7EKMONM8KlFcC+UkeuqNGgoy+PUg8hh1dlrHyfB
XWdoG4JqAVCqgJt4+HwORopCyaMinkx1ZemSNx1XtDoc3Gs5hteJLaqRMB6ebMmY
j//cPJ45wQ9CDJDgZRpOjCzBqvz3OTpcjmll0mmZn4wrjE8UwxqotwQ7c4KJPEo6
dKRLss63EaCZFHLpydnEH1AiLyNvl1fZpOrvLuQUuEfFvPc+W1L3rmlK6t9rdnRP
R70PKjIoYGvtDneE8+Wa4xV/FDO57KV+apmgpRj/HdLpDYvUZHlhD1G7SQqUBxua
pvT6lP3G0B+UuCkzyiYQHh3bQxd2RUtQKwh/UGymcWJXENEoIEFcn0cdkIsdFhXL
1qvduudYpy0quhEzoZ13IV74lOCghjip1CRcMSZLee1c1OR0k3OnCQk+rha/FZlu
dasYMtGVtm0r+pW0vZel89jBTruwuZJqaycrwDcXwu01tIalRz6lNfHC3oxpkWS0
+uLziyGW/wvoloqetuvLNF0bp6DZzpIvZVPrEt6Rr2CrlS1tUQ6WFw6m9toWKd15
YCdd6RyJPiZ0QE/6iWwgL9cVJGmQSt2ZN41gXn564LmlgkIgyg1QGb0p1kqMT8qj
3w42edJ5sS7Mqmgxcuy8WJXUhJIw8GuIN0r9IKcnUdoyqnNEjomO6fibKw0dpz/f
Pxi8zk4NKFWDCmT5wx9h949b7iQwgqnsSCqyM79SZ/hJSn8QKdMOJWYxqg4B0AGN
7JZUUA0OrKqiW3iQFJ4rJwMCIZqBub3G34dFI1W9Yolw2P0k/QvboXxqYwOnTbIp
2rS+3cT66NQRKFJf1Gm4PGW3f2lgETb+8kE3Tew9vXCwBJMc6w6BDA5/xWXFlFp8
dXYHh+sACVdhwmiiQzk3m8T1CQivCKi0vMSsvW9NSi1Oe+96M/Ypu6DYcqShta3G
ZaAdqk2cwaAwDYSpRnONoUHEh5Y7BgnvX96ot/0BnZ5aTdll3fmV8rXyIUBz0uI1
W5qfa3CFXI7HFGBmsjHmhE6GHMiuF4tkLVJLRX77p1KUDHwhdsT1ST0QIvFr6tvn
Jo35UOhOmKfWF7GiwPb/BAo+dokH9eMY+V1+GPiNXnnc0EBCm6XcXS7IcKKaNuUk
m+Hp/Acn463o/LjEQdtMM/YORUuOPIHfn+RQvAzJ6w3MsI+gqtQmMHrMLPi9sn7d
zAAdaFe+7gycjP5UaHk2kQ0BU2W5yWmQhGSDZtYbl1nk2+21FNy1ZfgsDACEHZd+
UpjJgUoWadP/RjZabXkiibBFFY8ULHtiKbu52EPVy7V+0QjmO2299UVRP5fzdsQ0
mtHjcS6CzAzNrIiYBakoXz23gN0kvakHYVPWL0ggJSMIrHtHe1yreMGItpcLsngI
cxjvx4jdJqWSd0fdVqH804/gbg1xuMtEHl7pX3y95W2TMkIMu27vWOZ5ayQ/LKpr
+ecga1H48QupY0LIOw9YSKBCPz1jvLsKo7/XTlu8JW49MECZN8VW0vrtGyITev36
EOd9X68UcqL3cR5ntkcpKABfTxyHj1Uz9IIP+zCmK8xFPypUADaOBcgrhfOd8CHn
oMLSBVAPbmStZmagw+O9AQ==
`pragma protect end_protected
