// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
COnZwcJsaNCWQG9q68aXg78vym35jXBU9clRyIb7O2sm2Ax1av2i4+10yocsMyX6
RDlDX3s2JOQSPJGLvIKtQEmw9uEuaPmj7Gg1PAn6pVXbBMEsq2cVMyNWOtntOK+5
l+IxJT0WUpwHqZ0yV07WJXh0zlp/OskZYqlNASYxnDY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16928)
hQTEj90yB8IXfiP2UWf5bBIDh6evZ3Gjx2c+ZU7MsE3juaY3KAUq23gXjXCiYRDT
ox7jQVHOIOzsm2MGnctUVlCDV6QOjplt3u3LIQVz6fU5xWWcLuNJfrks8+kNHtmJ
yNpWyDe3XiMOTV0vf2kpMEqaQ4RQCesahPbMktpbgwggyU3NLcHcC7jOsLRIBri5
Bsa5LqBOjg5FiUo1kXpL4Qb6igCtFTkAO5cBnKMEHTSgolLw+XLE55azfUagk9DB
2unzoEL6bmqXlflbFzcaF5ECvnsOYZfLP7uOpHSJmIzR2651pRilTwXdHvJNNkaw
tiPbdr8ZJaCIRhBmGYved0RGYFFdNle3oKHA65nGskD3cw9of+inHiPkJ0Ksk26S
YmzXnfjdt7sDaLwl0sGbjW2Ah72NiHYv2wsa6U0Qaehpu4g0R1xP4XmNufQqipsh
G4qYtYBVhJhlBDFWpObVW4R2E0R/ZpLCgE330XbKzfeQs0jDKB1XhT89sn2E67NK
PU0l035LmDG2qhMbsG1MbCDOK772xnXswEK9Sci+k3SU4iJkp8b6Wrm5H/EXQTnR
QqW3SZlvi/Q4J0M9v7OlLDxaGpDHN83uL0ybfc3sr5ykp8AeB1PJVlbtrTDAVl38
gQd8Oj4HB4vYz8KBqrVU3Y0EbqQoOdkSXiuWHl3TN4/VqVnSup2ENmsMmSNQLYwX
+hO3xfv8Pk9kbbOCxbMmy08rl1zaZaBBs8X1FUveYiVXG54QlOJUDb9IUe8gB3Gx
HK1lmoCPLRe/ZrVOguw5Pa2U7aKk8M1TKxKNzWLCv3eCCdKSPGwGa7+bflp9s7zT
OUWUXF/e3peH0EMia0Y3Q3Rpv6aQitv2iUjkCCMqUsyy5bes6XvqTNrTjrcrsv5r
N9ZHKcT9t3vhaMcEfyQcKW2JuswkqxMm6b92vXiskliv4mVYCbzc18vxvzZM28fo
EyR5ZR45jloDttuP1xqzUvxmsMGq1TgUrJwXHubqdbiOEs4gfD/VsQgcjmTOcFAp
TdN4ZfcdZourw8vskf+ZhUwHfn9fFu8PHkQEIkevpv0vQ2iy5qOYz0/XFy441Umv
7J7HmoIKiGBjCU1e3rJx6ZaefMKnkv77opXWzTWkynnBHRfnExETLS6E9QAqjnou
dWM/0lvjle29xW9B9z5WwnFrKCYhFFT+BgchsGVSGX8s9iMSgFElkHuj0qMshSL0
wzjG2euzWL6z66nrs3AbWRwBl1sCTMLeHXqxJhKc3xRZ+bjDhayd9OuLFEzINhuK
HncgSwE0PyfGMGhJObfFRNnngkE2vcuAgct1picXd7rFki+7vwQ2gRW3Fe197RQt
+GK7tG9GAU5PTuQo8JSdskXNvMsDKCzFNMbG4yZ7jU84mnmuk6cnUo81uP2C/OuC
NwytYeTznifQs/oD0itWA+qLBa9FWaOhOAXIMK9WB+hf4ik5HAn+4G0JJp94Cphv
RwP/9qCBLoo4Ov4GZCGK+SKN3PhzjGGKl3diZAXs2TfJkqrlQV6KFiA+y/ud6T1K
JUv6TYHC48Zfoz4uiq3gMgCnCIwUFjLHS149SVIls5OHrw3arIWoul8QpippMhKv
tvrscvSPoNqjjdQ65h6P/KecAuOV5EZb+supZq3WKuR6fbfBOwPqfeNJO81AQ0c5
0VtOkCKtI3hkbWtRMevuil0Ih+CqZPIzs56lB5M3ta16fnd/ymL5A8cf5DCrPDeH
aSCWwswjLwnPFra4MkssE7nIrvvZJNUulz+B0gp51kKvRQKwZJGUB53UctS1Hpop
n9g1iHmZjCr4Upx3VfDM48AWjsN4Aqi791j6aM+a8rRqkrJNOnWUJfe3IVnbLmof
ry1Krc3cc4tiIMl4JIkE7XuDiM/0I9YH7vmdvabZWLlMRa2tnP/nuLJtuF/flvyw
3ily6mETUEgzdZvN/wN6hsVtZM9aAwSrqoHhcY1mJWdvAxTojNkzU31xNwcy3euL
eJpNGTv2gY+VK4HISw9qE55cDI2Y+bNEQVjWhbiZr/E1COc73FyY5boZdF4ypfdu
rzsmxVR9Yh4yYLmN5BHiOEAbf5D0iMeTSCERdMLYetDasDKI6jG705t6FYJzAdKR
mNbVrWTUdzqOzMgkkoTYLQ5Y6BeevYU971QXGm9iMxil7sh3damoeK8GJ1xHnlg0
Ivzk7cFaaWNdfIssVxi5FUu/Q+A63aqwXz66nDjBJqJkx9h2vUzJdNlppkste/mO
lX5DEiOlTxoYDmHkzlRnDaqeBAVp/cRsW3xPMD3oObxoHH2Z/oIfF0etXOI483iA
YnJFKONJo7DUD/3wX1MghYBR44okqiMITMbz9tGuoPfbDHeicJyswWtlbbLOga6f
lseI/9wj5LIy6lmkoH2N61OwRy4Sl202OlekQPXSWQegaJVBUvbCCZfFbT8A75K6
6Tlk3mdIl5XAQM7Kd2ge87+0VQMRuW+7u8QcbfmG1zGpz19VbgxAgQF8chFZrTC/
flU1Usy1O/VR/6lNopZI76IJDSur9EF9MpMRyhclWV9l/ZZiQswKHtrCPOJx3LuO
ggWzWvcPqbonHoDsqW1MQhWuWkPnnnqNU4+acE6wcqXwM3NbBxL9E35NrFF7SO1e
Ef5ln8vdghqKR0z341LS+y03cKLSec5KGFYlRAgC4RUx9OAOebGtdDSnagdTvQSG
RQg1x3lDexiuYcQYyKkNwoZvIp1nIKtqWuI2XT1gf1n6qPdPk/mWV7zyqT8vAQSM
ejegkLm7a1crm6xgqbpOmpztjRPAkJMj8nE4g+ZzlZhI1gzxa/a6zSx63V+F2kVs
X22f4FCX0/nsaMkVTQ4SnFO+HTmwGS/bzIHbvQmn5XHu0GcQslHC9KuxQV0gy8LT
dUgDAqU+l3lsmHFVhLyVlanDPvOQHBEqJrF8F7CSMiU64UdtlpvC2fVWj+WJJzzu
c8mTNSW/e2UbLyWYHMo8LBk34eYpmC5FLVVdr8521YZKsJH0R43UuODJXgxn5DHq
4gu9bEXBjaimyxbNDmFDgD2clyT9/LR+ap9aMEnBqC/M9BCmu5UsjnkTv8rN+3kZ
txJorvCSHPp9xyRGTsOw4UDb4NeHtZ8YzRMow3N86ZgbwjuFml8c3+nQYjlV5Y+z
/+IxkP5qu4r8w37FIb2C0i7eS593MBKmE8fuLTU03/SVRnSjKkVWO7+RBctg7lSC
CLAa/Kcxkn1Qzdro5UHet59KFW+7y2p4oyFMkTcMukj42wOhQmDoP8xkEAMJFu5R
rD9DydlGjv3fe21jhpnbXBh9pAeHRoXxlZdnTk/JWySjgCYHpdBcNIT2E0H7wUWF
cPFDCmAG0jwsqmC0yRpKlP9ovMSC3jVc5YfCrh9oah67qk3c7Myt9k36PjobzoCZ
uwvoecBpTxh7wERIWCoBIV9Ou3z+4ed2SfzVCzcqYecGYlZJViUSAvwR85+GM3+r
smr5QZDkvaWhX/43dkcrZDEaTJ+tlq+fEQIf9JKje1WYPnJuhxt+P0NZzk8awnHD
rTTxj/2oNtG75wZq5dxRoHjbU2Zr6ijlRpmZd818+hp5vRdfAetLqXJsQnSQ4f9z
wZN/UMlE9j7gQ4t9m3q6WtVA7iS/+3h71rddm/8coTI9uAnwOn3RstVe4YWTOkKL
BeQK6c5m06zXNOdo9GnpPLrobNClZNyKHqFsuD5DjFNRXhqKXBlZTG0xkXoStw4E
b6nbWg2r32KGLjwS/taTJK3WBgg+wwI5Wt3JR3697gB93pJINwlGs75Nzx2bonyO
wTvIPJ3fRMF5RUqfZkywonuqVd55DT3gE++sJoov+bc8G8Z3uO8+6BCtp/QPyYOj
mrhsYrSKANJ8Nkgd2ofVhuDAQDSg7/GE6R9aLUEBN4b54PkntnLYMWyV7kF89v/r
YythEB+uTZ9/eDzD/ETXR4xLXXsc9EbFIZioMDHTrMx6UE+fO/UfjaKGne83EnGz
DuNMxLErf1uCBF2h+jmgUnhxoDxDyb/wZXG+55c7pPJAOT/o6Ru2T1ak6conJ7L6
gIWsl9xiTMu/2aYwVnOrC6Pu+eHRPBt3C6P/Jeqy/XbiWLgHiEgFyRpy8A/65ynG
nZiZ6hZj2irPmTNS3vXrrf/1QDMraUqPV5oCj+gh6BFJW3kq4iNWPBqRQFRt3wGv
Zn2vNfVXETv9z8BDowUv3vhTfkbWkpxgOHfhEBI3OwJnSrgnC2Th7tNDZS7aQmw/
vUrSU/Ze9ymrOo+ymhdzkVYksF002bA1v8ZvmViQdpo/TGbi6xL3jA0INUDT+2Qd
4chgpPFZ8OYei0pFYty0M0WsDPB8Vqu5lkVz/rLLPWDvXXX34/F2HliLHruYosuh
yOL0o4UAeGuHqHOZawNaAqSSoqz3EG9MtJwRnZ09Hlr2dJPUsrFOxEmNCSAoT3Hh
SHuNbtl7rxTdt+HHpY1Q22H8aOeoNeI/nxGmOO6Knu1rJeQ0VmfXucWuNhIeZhTx
L5NPAR11G1UnH4ddA5nDkE36FwcgOYJTOd/iVoJMZvppvR2iU484fccs0JCde9Nc
S2KeRgecbYfpQh1Zl9PxQjA8nYTeL2jKB8gzRNoeQ4NqTOZ/gMb5DS/hkPS+Ov/P
Vcv4hhBeuhZyuUuUoOgmKPKuoBvn6S0JCgxpkGm/m8jqpHDtjjhNGb2v/lsBqQCY
gxXl6vRHiwcvc5DdxrmqDrPu4/C3juKHlpqhTLLOtMZ8HMaI4nQtyAoOyz5Ml4GM
ba1P2ziRAy+AUbOlEst7nHzV4JcIFfd2g6vuvGq8uAXzIgw+eJl2PuhICsE4F50k
WldrgJaBVBE+lc8dU/kNosKkyilaVKCpp3Hs0z7sYOWTT1CzlDJm5UFdSSrarA/h
R9YLlmQXaTD0Xx1xo6RZOmlHSR0ux2vAjUeAeWXlZUOBWS6wISxsjQcSnq2HEp7T
831SRCI16MFkW0ZcGzkxE4M98vjQto1bJcsw/Ot0nOAcymPdI2i6loxgzxFs83bz
dGYKwnV9FCzwjUwq3xL+uLU89xitYOFLhaCxZzWzlK5QGwCW+74z4l2tUY5tLzgL
l1tJuwi9M89+nwmhmK6zPglc9xeII68rLiJQ4QY6MRX4BkXkkz5aecggefvAGcLj
hbKiCBcuxcT/6ZEDjiBDIPsX9kbWFEsqdzADmQ/6ZZ3o689FyJzFRiGuBsH9zDOp
dZvLFhsxt4W+4CV+J+hiDWvNXHoCxc9asndvka0etT5B4Srl22FpzBhhSQG4VZtc
dXm/vcaKCNT0TMRGKGiVy1przVWe2aEZzmmD3ah/XPO0jvC/eMKT5o/186pUwF16
OKXlc5VJp4HOcsHgqouWPLnmg0b8DtMvpRGSn9p3yQwwB0RoCK6LYj+bosuQ4pbU
t31PDtwMwSb5E4apSv8pCh7P9RgUxbQT/qrTysUCIuu67dhRcIr68VqFrAJnOyWS
ycb2cUjYLuWJmmot+nxbaSVwB/YSAmlxEtSO1V1AgaYPdqL1OrHnCRkJ931KaJLj
N8PEER6jfPJmASS4IWzCfHt2Ol1fneJ0RnfrN1e/7/t5BNwzMPQw3C+d9vCRITml
XJo+cjV30eNwlIwIHdT35sgOSmt13mkAH+ZQhzobgRwh7nzWjbiLRr6A4mLhI3uh
Acom+goL4rO+CDyRu99L//LpZ+dN/hMKc8Ie1iIoWP192807q6s1VIWWgkHO89Ch
5w3LAbPIG9Z4bxDMkjCRbP5TIdAO91eZqH5Dt+kdRmC7U1zoe8+B+ZFeKzCHBFIy
WTccYcsAkqy8kbJ3gE7QdiWX/Dq2DJ+TnhGML11cUeR3/LGcCXZb14OC5L8g/+B4
iQc6F/RcJDWxbvVi0mjx7QtmBO4vAW7bsI4yJIWhhjRoktlRXM2sU3nvu/IFZ5tR
eQZjlZDMut2WUwYvzJkOj5zGwe9X36O14gKheYww3PsyPwxDEVOPx79x6fbD9W87
ZjxWJb1yKH8XBIBXQQmOTeqRV4KIxbNKaHU4wypft2ho3bR6NDv5OHE1zBahPytN
n5M7RDrUKY6B6ir7iPDzGbxrownWN1guN/3iLrsgvN1+Jl4gFlTAtoQfINW2T9Jd
vhtyR0qYRiDyi/VPCtd+7YnkVoGdJHtuRlzc2C8kIe48tyStsyPHyyQblLL2OjN9
hEYnowYy91JPrEDzVQwTOj2k7yzZDuZunIfqiUb/tlCdqOncayzgzEuSKEbP4Bhs
KMrSTF2vwZ0p/YnGckunE25Q1N3RxcjzklHPgKI1buH0pxtXr0yEcPYTxytoFUjN
Yl6iDogoo674fecx7956yufeMV8/gjtGrfxcB81XMvq5Og1+LQzaBQDsZCyS1FoN
UebmIZNUBYpcYs7i3Ybk+kqoXQ1WCTXOr38vPuSyh+uYapd80wnfoYjXnCzE3kZ8
hq0jQu5uGzq+2Iv8fCp6LX9hFBtSqM5zSyXsUbfqIPVY/XAEqnNx/rkCE3p04ZZM
GVOWdkjnU3ptTkHpuw9yEOzJ4hTwu4LfGz7apkaxLrVh5qFq0NkSCVQTly7fNNu/
gA1uU6rL+lk6UQkJofN3kkpwXHpR6XsdpR4SKBhe73cHyMzyk0HIzY+xU9x639jG
+GeDHo2YGRHSebNVz3IvNjtYbD21Mv4CaV5Rfxn/VzvWcA/d8riuWEGKfSHasIFO
hi+VBAnrTvRwyJgxVX/Ch6RMclde9nLsZFxKIoEMdnjU/inOVPPtTIHrTRe8eIk+
ieyjyaCNkOQcuD8mvr7RxEimPHbmj3fxBRmzXL8S1EY4VCJPIKtqyAhYHFeGzVcv
xwFR0wCjsVNH14eW99zEi1qZvBtiSfpmYvYZnuIsRlYZ6+lkVUL0ifQyxZKVfFsB
RmnbQZsd6AJ3XVp6xuZ0y0AtnHRELw+ChI6L9AQpKbOXUXvG1CRucJqBZ/ykLgI1
tFnlCXJi1nqH1T0O/RJfNNUacMtzgn+ZTMnHWripa+wboJWkK9LGsR4VYJypbx9f
pECpFtONHjDJR/DERU6b2ZMZQSaEfVe6yF1x89+nWRrwhTSDOiIW1LT8vDc5IplQ
VTUE6cvuIGvEqXebVfha16RiCnGGJbm4OkwAh9JKcLc4DiPdEsEt/pA0SwIuDURb
aFE844acFO32Z73ppPNEIDYsrfO/UfYLNTlCU2JmraVTC+w63QTXy6/l/TT/lc5k
AWmqokiFG8Otw9PpL5H2PqZR0xPeEQe9gLJ8Dh9Ss/NNWKH958+CJUjkLSOfM/23
+5jF5szvbwLc2jDxRou9CGj2ytfRVvjMsfb2ISBS/4vApAszRi9UlSPJy4oI1toh
1Ry9NLhlIVcnBN1dXWhYPqihF1lxJ2lbL23SpTmyZyxVaSoKEqrUeZhm+FWit+W8
Z716axRHkCxnUD7htWkkZg5TBHsYTWClqfM7ZlBkmZkbFfo8/fc61rman5pCjyH7
KRgE1wKLGP8uDNqcC0vPUIGYxZrzqFJT8DvOqAK401fMoMBw5/YVqN550IhrAYDk
fCivqaxxACM1VTBmAisHFxSrAqqKl3DcP3tvpGxdsQGpyYOBdTeJBFQEEojfoklh
SdNlkfFtH+Z2eA+BgUDtCvd3YoyjUyoWYGkDFqNvHmMpFUQuMbLDiJ0bvBH2lLQ4
mZk6O8rKo7zUMkdnKizzaQxAUnfJiaManuSyNAcF+wpVH1RnlRCZNB+cpOGc1SLE
8twNabdPZlePEwdmDXAEGqgHQjWdWImV58lr7evfoidEPz7caGEd0u14ebYjUstP
FQx+0yMMO0ikioiK6IBPvJr9puyRj+VgDwhx6kvlqcuTgw06jwjdU/xka2LhoKFO
2fENIhVt46xRcPfVZKjDWHxIU0DwFz0FgnHkP9HEHr+Xy/NcrX0eryJGvX9RKhHG
rH3y+umEBPNijEiVl2laxkdRm16v0fTrhqx2zcSmPBoFXL7zQVXdVfWbRnbMErrL
uzZnP37//eOipyMSD/lGDr2WPuo6Een1P48mVKlH4pENuD62MAF4kokJ9tVudqCL
YEckm419CYCnXCUJA7Qs21JQVlhfD4a7HDMOTCA932EW/P2QKPfmxckHKfo9aMYV
ZtSZrSOTzjRZbbQd2pw/xqWtUCtE+3YJ+3zQPZy+mzfGogB5bCeWcdfhFSiAyIGW
uILhqZX11foTstlf5Nmp/N1DT2qyf62aMUeP8w9r6Yq6oynrEKioFcv95t60GGL0
sXosUfcDIOQjiiTSZX/3yUd9UAq8Cm3ejnwwn7UVA2R4uYycU9eH7u/WHT/IiONw
k9ohtP+1eINLPvSpcyq1Sc3eznhivtfFwCdrif2talxlQCw3L6blUaJQAfHIRp4A
4M6Le39P2FOxchEKoK4JBl0ZVECG1tBGZkakVNRlAwNv8i16HgtmketrWTOwujal
nuH0vztIkRRCRuLLVhgzMX8nFotgmlMlIzmRqPWuJuLf4PNa/mfi0kG+GSvWcMLZ
WitQN9kaoBFlMhL4vVJ7NEGHxeBg/QguIWxE+6H8z/Emryv82YrvnZMXUCG1BKY5
uQ1xdfIa94lWefLhVU8dbpMy/sgpq13jufHuaggEQ00vwhOdRwnZbtDaVwhDPcQM
mJQMDM0vg0db8KtWeVQP33fl7bBlCqwjf7OhoVZqKieE3e0VyUfVpI41w6H/Cube
RHUrRWT8DorY+xL7drMD2ePd5ksnyknqE2Pik1EqRSOmTxXhZpd1sQeQutIiUEhO
yX8F6ckGDLcw/GKJE7YeXQgMIuHg6yLWgO2RoUxehJP701j0rqWCac4XTRVkrHuh
z8WLctcGTghKC7bbexZg633PECGfPFdqia/vKcekye9rIasUrsqZdLBl1h7j2Dj6
fPApMBKsB0PKTdWSABbZ+SsmVTNzsRlo5PkeNzYE4N1F7RzyKjZQ6J+Ic0KmqDZ9
w4Zyfms55jowW17PGisTw86guCMGkYrou2B2ZgOIa/7CBUD30kyNvrYtZ8toAe0U
t7zXdDFbQAVeTcPpDCruGLrTWojz5JxK264Q7T7cKC+wrV3OD2gJFvmW5vN35XP+
6S5v+oCFIFyvxUCAzUNLeOIviQQzODL+xV87ekZ+qfEN6SlbM3Tlq1cMr3S6tWPt
DI+aSmoRLpvGW+EyknShvJvYWtbxDuK+T3qqHIk8LQD65z3MzJy/kLtj3E2tCnL5
rpBJX6B6mUw7O3c6ppQQzomxdCfh+wK8escbHv6SVvDPC4R9IOEEyaPOh75XGGFS
MC+xF/iRh3DgMM0ni5I6lQZ2lf6U38x2ju2DuWU1vJ8VVmfU9ce20rEd6A406J1+
zWf2IGkCJaIXJLedxORJ5Dt4ANr1SOmpEcKJyKVd3RIlhmWhnOrwlCGNPM8WldWK
c57VXdwK4g5trs83UWU6PcyKjUQOhV10vaU5QfCb6hg5G8U7yoPCWs4UxdRBHEVQ
bMME2YD7QP0wXtbHod46duuR+B5mk0r3uNhgB0td2LuMrx6/o9hosxi7CSahJ+6x
PyE/WITTbDKfkTZdoBVOYUsEC725dkC5Q42zMYOVcrimO3pq5mmqHktPPrCaZ7AT
aWp0zzzr5vKsg1HNS3Hs/pBSvH1fHY3w8575gVQiI7D146OrvT6ME+HdsmlDRLLb
5qtSCkWe4IrOvsyisTl3dzO7LlsjXf19H4Iij4fRgU0vTYoW9RE50eLD1qfOwxyA
dH7WLMFAIIX17IsYOrD7FUkEIlRPJ3Xg5DIN6r1a1U2Tudz3ufoknAqBG5zb6hSu
UMIAlqh7ztS++1GoZEUcybGhu+azOiKDKWE9AOtMqfW46c/18P6/iW4Nfz9+voDq
4A+H8NPveJB8uHdcVbKLizlAw9ui8t4FXPKEf34e8Z+oIRXd++rhCO6AhUzcDjXo
qoF9EahXL2UelORFWJVifwDtJHVMmyWQxqQkbiQnEkKSbngLdeSSzhp+9m/i8l1/
faIjYshS6tQywH462nIPCXQKoaofcYKvbGV3locVo8C2KLoUIuwvKBLyL5qwKv0x
gVWZkHKjjr7FMJHINEoLsMvZmMdvZkyew/wL10B2uwoPvD0j4/LWrMXEjvWqZ9aN
pRrTHFmott9Fl1p2BiHIl2fWiFrBXSZ83H6B1NOh0kd4KUfpfM8QmmVQw0CuS7RY
OyXQx1PNczcvLaJFE0+B1s6JlN6N+Y5Vsec4uVRuBYkK16Fsyy0xwgreyebV1Hw5
xryKztDd1pdaJ54N59ejNiwm9KpgshhqrsE+xJsgmPVIGCfwJtalGz166pHwLoFY
X/2lWVrav7PnhM/0YfDLcjohTg27GxgMwQS89hbgnxD2f3vYAZNQ0SIPs9PEvTj7
IjcL2zUCs4Z0EVqLidrgVEe1Azz5OMerLZlHGHZYjM1mM3I0Ob9s56MpN+laDKfN
eUPuHlPNDNRBm1bR/RzNDoIMeKVIbCBP1PfI76geLQFMz1Gkwajt4YU8NawMBq3d
eNQrOm3Scq1OdPlHqIvrWips4O/OCuEi3hFUEUO8u3Apk3x/GeDgw/QCosBOSAiF
QL6NAddArd1pVjIcmOmnwpl1+SmlEJmAQ8MdzGKZnG9mNda6bBIgP9kOl1aKjJGQ
AkoTS9lEBwfuMuTQr2zSCM4FE+IPnP8vT6SffVaLRWlvRP/OF+RxHFSN4P72Dswl
eiRU36YdE9rDM7WU9MzYXqyt0tVg4ulnHwl02VUEPqMcVxgOizPlFnBujzAzhuMB
kPqL1n5QCIHv95qLhX5VqbnBXLYXp8Rlcc+vCA5eABQ1CmBoDu0tnPkJ6E8NJwAt
xnBForgRCrT5wdGOC/Mf53O9RCPHl+buVk7kfSHKkfr7JfmbH794vMG4xpHotKnP
rcojW7IXQDbqYdEnsNC6P3+QzuIKmHQ334VQZNC7rrdZLoWb4+Osxd5LSYdx4/AA
fhwJicZR+QFzE0GzK3Gq/JCoNz5lEWIJZT67/wNADax20ok9MXy9FIDEBvfYUXeM
nNy5cbVcjrYiMOUMLNiNN4KXci/Pq+kOGZDhjhCO6VY6OPqzPEGVpNIXh1rmk7pf
meqHzjuZ2lgse1ED8pf/lSbqTnimPLpGLLgqPSZCZjZN2+oPu8zYoQ5skUQb9HF0
1ERfMotAZi7hD2vFuGDPVqpQgn/kj//xOi2GS3Q727CDjvji/PyIA6nNHGkVFlNB
b6g6dO1GHWHnL3Xy+nzHPcudSZKkrYI/ZICgKZM0Pc558U2kUkEFv3q5CPDCJyxG
pKJTzm5ApmcfHb6PBo/EYQ9V+W/kxISw4HCCVgLOb/d0DuD2QfxBeUlt/+SFudPC
cBH0kzIfYrdJ3P/G7Mt2auOGyIcLAo5Vi1V+//GSX1cONLk0Pnn5GdpWpUMiYYDc
FzXw7ElHz5gpcENsAdLTgdMf1Hwk3/hkueZtzLKHavGTZfIUgzq54zOwEJSHpL46
OQ4Fzt5C4f/Bix4AnyPYxVpjlBCS+dbAlG4aebEKjH7Km+1FvcXej2R0fTNIaNri
x/G5fqOF7zq5QQAwN825t6e9Xt6QKycSynvfX+yQHQe0ZaEKotjRfTkvPn8fpYzw
jNWIwUqGNImMkM6YeVWHbDK9flWNyVP7dt6Xvr5OqiIz9DS+iPLKOIkMbrQUQ7P+
Dl9KziU+ompft9RYE/PlEDyhUezRg/8djTJmorvdUlHIbydxyGuhmApVRxqGQl+Y
kiWcNcHl75N8QVCvqDM/C2eb89PXED7fhhmUtY3BgYS1cv6TihqmY9ZL30lyTW5X
39kdsIQxtdzFpEE5uzdoyxgPUB1k9f1RDXKKc6fKLxY3vVNVu+LKRqDh1TinBs8n
lDTZpBo+Zn5NkVmF28C+SO7UuQciujletSIXRF1osKCZuP6tdbwKL8qAEwfJXAjM
r4YyeS9gT8QcB+g261j7HV9s0iDROi/p1i6Wh8njZ3kECtZtqAbxdzgidLIxhGlY
3zVazyOuhH2Lkl1lefvV/VEFmqIzMRcjduYhuwVig0ZhITaPKSQMuDDUHvZ7uiFA
4Qm9ndzjuj4ZiNrGnVwCpKX23DN+GQtEak4ZiN9VeYjQ4Vgd2r6/BJPuF8/0uqXL
9ALkhejBXQFwgrJ5FujB6d2RP1w6QvF75YRJ0LIpYzqU3pK6hH36w4QhsSy+CdaT
ehTz/tk8CUYPmywTNrvsH6uleAqXJZ7bELbTR5BfYh+S96snJwtJi4RmHI/GQ2cC
de08RJQ76mLcQq557Sx42fFq1LWvhVEeY8TBhsVOuDWRw2qxqbTm/BmT5yYnBUye
F6TaSRKyvHj5lVE+9XsiXiaHObMFWo65r2r57EhSl5E/xJIHhfheaaQeyf9rLutR
m/Yta7f1MJZcejO7uFWooLhUDwVtnqYLh05GUoI0j455Khgt+YzBIMhhObC0DveE
pHQMfpkkq8gVzKoKfxxmeUKgI9xt6o+Pt7qQ3Cs1GC8YF+3KbBM2Tal6dN8nbvHO
cp2bGnSl9ldcLgax/BjScPocZLsodgxzpCGrojE/Gtk89RntcEDJpNoUYZShBIcS
+RmCM7wdqdabKNraSnrv5i/4aBub1dyYTli4rgYa/JIC6DSzEaKi5DLdT1zZXShe
eDVteFDKy0CeoN8EtSnA5Ca5BXmOn61XACl59R0Ft19cEsc2/w0wkEkNeIEun8zH
Pj2v/g1n/VyZRBvUUQPO/wh4Xw8Pzz7g+I8yBuraaos96cMSxL2bvPqcPEOjuHe8
LsxOYyazy9MCmxI0gvOCyEAn3ChhsdWSyZPM9lbSK+52j+7ClOE4MDT4bQlUoLv2
fijs9JXmXBm3lIhT5Zf/z34oWHxUgzWYVjCDAAgSqXOTnXU5MNE4PU3EqBVs7Lgd
XoRyh40w7PVaFzRa4gzxaEIT1RyGSDS7duQq2hWV54boUhgP2ZbI2c3Wa15uQSOS
9UncizyHEZ+gNlqO9gBxPz9Vgqwq9xanfiUJwmSFGWZb8v/SCw4tbWVzftsvZ3qH
bf0IxQOmJihXiteAZlreu+dmnqtzFg51SYkYWx+jSx5M61NpCKNbqIePTezbPeoq
eqWb3EeZ642tJgAPp+RxgXLxLdvLqypWwUrlW9B6cJPSyPX1kmaA3Mz+GkLookEO
l4BOy8o3ntGUSfaF6bqLy/FP+DOh2eck4rxE5m0vo2tVBOSie/UPP5APITXUzsen
1/JvicZxW32/ge7PKVQVTxQfQO9QFYhOpt0Wm86sdLHTsSyG1HA1gP98TBP00UJX
aSA0awDlaVb1BYzcs9ginp234aESvFIWY7e1mPU+mUQepfw1vFd7szqQmK3P1qne
lPC6pKgujLnLgJd7rERD/UfeQZjLIuYWEWOvrxgVnY/pAxw2m94BAc9C7SqAcsSM
4OM3X8JxwY1i1aQY4ZtHDpBNZg+ZE27y7gO9SJTfCwASVuLTobpSC5a6tRTmWFQN
3WK6Z/93RWkEbXRTkIRht2as2Mag8gKv0hRD1RsTtkFLYXaQbMYmuM0t3CmiEfoc
EdIUF/8XvdEdqfRYtVW4FwY3q1nBGzguiJmy60/7+SpHTf+ht28FyF+4f3eC0Xae
rIKALR9T8ao60ZlM1fO+ujxxSRVpRSLOeFKFDqZQ4WUFdVqozfdyTqCpZYpr/dke
uOnBIhBwvKx7Bzvyon/hcvcGXDcioIqIKydQLv4Vv+O2+mNFmKlmM0ljphM4um05
4r/4VFLZCIB1VKkid6kO77v9Sl/wnjPeRsjGqmOjgGNVDlWjyUVWWiBy70SXlvgp
AsWApMWl4v1jsIQA6ZiDUof92zOHq2MROSVe+L8qGpIqC80UahjwOtsGL3F9GiRl
32tJw9ajfeV0odjQExeFrP7V/LUmjvJD1YzyS9IIdIaMQObYiYmdqlj8pbtyw9o4
O1j+XrVCbva68A2M7xws1Qh9ZoV/QVEl0hphGGO2r7S1EvDvwnzAYyM8/lw4J24M
NKji00dBWCpM+PyKOcSPw/Ec9twvHkqEO+1pmdhsaEw+8tRv9227IQXwnKm7wUQB
jqMBPIBIzmFxntQX1AUjleuvhPHLiCLX41yDWsilod7OcB+2Ht2Sux9OJvq5YG2I
WHzyVz11WEy6bp9+c6pGhEcNbQtEjUFU3jJvAqS9Y0GO27yAOkhw/E78Ai9bHejT
Lq51MWnvgEFsFCaoawTBS0VS+FP6Gg5zL7kGWV4t2GfvwKVmiYYzQUUvScRfKnnH
XIeC1LJ004S8kKGl6dGergVMwfA7NT97aL++9mWfXj+5gjB8wjbI2iU+jBbEYy1t
OgDNOZPG4wQqa9dQl22N7+1UWu3srnHwadcMaaSX9W6Q7uXULqpKuWE+Y0eVVE9u
Ejgv5tIuqqDad/xFHVpvyDT2j148jtmcEAI4Gclr8bGqKx+xlctsSGC0f+DFdV1v
/TR/1vtrWSat5ds6YEI01eQgF9t5+03BqYKneXlW+HgWgnHs3UDaRJ1gPJFhhuUi
anyELJfiPwAwZk35Zk9ZQ4xnqVcfn97tDSdzOHz9uB8JeCGfApF6NG+XvfGYCp5H
yB4s0TLhoq9FzK4sSlmqxjuid5w5+NPJXAHK+UoC6/uHG6mf3p75/oqV1WU7SFru
ccVwPQILAisBXRtgiFVe/DB1bUHwgtAmCpB4hQeqvHmToPgmMe2OaKwvqxroGmEs
tMFJJABH5v989Tm3269QaYe1fMJ00nRf/XI21qtCr9X88MKrctpOx/h+sFFDtoEl
Z/cgsb+02+ZGPlyRcTQj6bbIcOOsjqyGafXGh5Zruu71lXfO1RNdmV57fGfS2lKz
SzhecUUjuCLZsoduVGqW0Ymo3EZ/o4A5XvxYT0P+RkNpay2x/Nj1zJLhYn2P3FlJ
IhqEbbwD7UUTkUkCbSs9p/Wl1TmTrU3w5hrOIkE7U07CdNXcbq8YF6ptLuvWyII6
8NXn4m8Rk9fgaXIPp2rJrC48aNLeEatcnbPeN7L48WaEdMIk5cMIVzCdP9d1Lk6b
vrorZ7ZXLNR+IZxWFDYCEwvU8Kie7Zbm1uOFiPAWZ6oi176v51XDLAhTfbEKo5oE
Xx4/sZB/HWHlXgpjc4lp8cdWczRBo+rJIdAVSZZLKx9qaiXyNXcbKaOEVg1MjkCC
jrf4mYEMPBYu3CaSbJ1yCU47vkoiMaiPQ0GqMlhsSX2cK2WJB02MiMWUKBv26v5F
Gcin39usRKDebxq8VEmK+GyukScWOUInYQsMQQhwVsDfmH+rnDOrm/bt9ODAI6lr
Y42DZEZdUg5b7pmD0INPOSaSotvxODPC6spr7WSIwIdz+wXhLrq70z0SDnjE6G7Q
4wjf9ukhNy2RK8fBfTpB81wV19Ogx9FyCZhNXZ7hlWIuGIoGYVnKO+rWq9ppIkE+
ouzrPw3CeS4IdAWIBAZenZ2Ic9Nrk7CuoQoa/AwDXIFiMYPFxRVyowx1UlfP0Jen
u7pzRp41nf6mDOqqgU7FT8KZQt6JE8wGH+RN0+pPyuC7EifHV+aU5jFC3z6/qHCP
eTstJdXArnZEXqImRHHY/jcXAcowQiuq+VgaEm8QETOTiIDjnIAdW392d1rw6IQB
fwl8OVRSsOGQuw2x5o8wDnkrm9BCCK6TobazEf5/NJKz1nh5q2/JAaF1/hQ1lEQ8
VIno19fZphczGI3nsO6tFYy9rbKYgEGwv5oS9ofaq4pTc9JV0X5UAPzfEbDcoKx1
WM7X+CJFHl45ccjYoChrN+1PWEHz6ta3ZBXh9n+THHEiJd0q5WgPtLA7n1tQIAXj
Kj5xaYd6XR0A6s65Oas+VAgKOCk7e0JfrVD3RNCIA9ZDDdXPaXDnHGtx482Dh3iD
BlKxVNNFvc/MB6GJqywY8mgDXdZ5eDtuexmpf0vcoPYS/tPJi1rDo/2Lt0uNIY+m
w9I1H6XFc0OjT7qHLoS4xE289ra1nY0SJ8pvjar//02LNgJQFaLYOngBSZXr3TvA
pH/P7R36Ti1W0NNMKiytj9L/77baJPxjsMEGlPWdaYCoNnXVVF6Hfna2/8BjctyE
aMOV2pTOwSOgbEJ+tolMVcdrgQOwYqZ71IV35NBTZ5/KGx/9/Irgv0atk4LgecpM
jQ+Ftj+PcVvhjt1c95DAczNC+qRaQEmJzWZ7+w81XjSfzVUr01IPQJfRpec1QMgE
beGlwDkDF3BcYqKse8g5pPUD57assipPdDR6STNQ4k09rUBf7mjVeBAMoBVMtXZ1
n+3PE+PxjGWESm8xHSH1EpVUyw+AOMf+fhy0AyTlQY/uDg+yOVKm04NdWdtyAt5S
Xm8zMlM5V80wXlTdSCMSkmOjcmmwJLJihvkbCLXZ9gZ3/oytkiC5m5u6z84tMgNd
6GusUc1SvZfHHFujN5GkjX2BCU6+avOMRciOq3ATNTWf2hnLzgMcxzKZlRk3LQsK
r3nB9xFfpTRtxtX29oPyXgSdBhSwG/CblIu6Sg3iyHegRHtrcd6ciIymlrskKUYl
/r01ISjyeCsRr+XN7bsg7EZCzxTI78ZCpHbWVVAL2G2kAVLlz7E/N8tZcqcMxa9g
xIUZjzXRDVkpEwJAJyOsXBRvpyV5pTg/wlsha2QF2rmQ/CqOUbj7XJvFcHwh1eQK
o9WKTvYDWm1+CKbXbY5CoWu3P4u2zDqFyHvdTckRixFHR0xkjPQiI1c9d4Pog+AW
+pApovIz1np9dkr8Gv/huF01lBdSLe7dkHpItrIrJQeYPoeh8m9WzbXrceRFDZ1i
5cnd120tTrwD66g5VBQAsz3ln0FOB+q3Ytq6cQWUImaQLRIA1RzDdVC57tx2zXB3
Zxu7TqPtYKIbGL/L9CBUEoiMCOA/0Nh5Whov+caCoki0c6lJprO/vlObAzhRPNiB
LOX82bT7hr+P859p80P8n4E7kHrWKAVxgaw+2h0L9ruoaiZa+m09XPzPXAbKfDTJ
MEznC/9q8Zwx36zaCm3I3rbf0v0I1CCv7gGWP6LDZeg/haHnJOjK6zf9AzFyoVhv
1GBveYZSU26K9ozeBjqVm9Fbyt1GRLaYaKzQk1OedlzYb1843omzMth/77aiJfeL
+y/gSATrd2HHYqtjd+UJjINuxS7GoyEzAq4i0z2AYaKXDJf4hHXNugRuJ2rYQg0a
JvujicbQb5JiOrZQEqxrOtQf8cxTVQ1FpcHe5SGnXseAsdaBajwBeZKCZK5RR1zK
e3/RRPowapgjDlZYPjNm4izsiStJXBhchnN2Ofi3xJy8H2eyf+VNrVYkA/8A4TUs
Jwdzk4lfxzKHN4FC+8ZGlL0NERM8vDsIPl9tC2oPOtmAblHzpUxhGqR1qJSy30NF
e0LHn109+/YhBX5/gqSXFafsTKTXkZl54gyQgwVA8nMrivzgYya5DphdSP/PzJ6l
g8RnI2NtAUmVSmT3nqSltRKKj+TyKJutExllUoia+DHYMcLozN8yMph5FVoNwwXp
BroZ1sfqx8Su0MokU+esFc3cWGBEJRdwfuF707gqjEnN0ImXLFSSOxkSt3fiNH3X
x2+jY5OlloDteLLgl6vQRjt+PQuGSUwEkbwYX8K9PUI5rH1jbbIFnqAD5T2Ysz3Q
qW0uKCIQik8JrO07MrqKv4jCbezWxqvq3phQZ5duqSyQTntTsgpQ3yA3M7mRCsbZ
TqBRlfHbH0r06u0D1vMYOTHxlzsk+rjpW+vxdikacgF/jPJWCJnJXNIgYhgebqgo
N2GzkZJbtKV2zkrUe900zC3JN0CD0sFLqKI4B724dofa+Fb6oECtwZeU2apVxIqz
7S5E5sgeuUzH4I9EkVvMs/7NTRS4353zzgPMaiRdBGYznCY2KWQx4GgM/qwSDCtY
yc6AGYBLpekaagbNW1D8tvInEzos4P9CLZ4/iIqjhgmAXJGcuik34g+vtGPJjLG0
yh1HKfLDA3pPtRFaMjwoPLbVMcXYhu942HF8rjL3gAYs0XfjiH7WTHjW9ZWHivU5
7Gdrzm0j+iipR1+NT6OkBb3vktdS2SeUiwQXb5gVtv4pWFdy0yec7l8AtGycaRbH
5FIzdE0QkkeGeRML1wfrS1Tdyl/f9ukQde8s5K6uG6Lwf68SFfGbsJl+3C3EKR1I
bi6RTBzcwFSpQKpTJukQ7Fl1+VkFJL2K2jhyutIoADjmGw/XsKDdm/2MSfo16hwi
sGYVZp7j2HWwFHRfTdZMjulyyDO55MFXjWUXrJ2LzO0AXGNXv6fXCHdwDDqXRcOd
MzQwzdOgQjFknhQpMXVMHwYNb53qh5hqx1skT+IbDH/jxIhMmpqTSBugXnCbc7sy
64/8ojh83qHTCwj4xJ1nf4KJyNsiC5iPOCCChm/Qlj679p1rFdlhoSXV/V3Eh1gL
nLRgo+pRt9vmzZj88bLksMFHB5lKy9X1JGL6ol6ltFwAkzyhDBcwih6j9yrzxIp+
n3hpf6NoR0Vdj4d9WjXsODZLZCG8VEO7hI69RroSF6WSOKPKSIqZ2vTATpOj36kF
nT/9J/1IRKqpLpNjpi1mopY6pzLhaUcP1VVB8mix2sbthNt/xHMDJTv4JSj2ryfo
y8MzNUpIDL/S8zfQ4AONWvf4NsUbnn1ujwRA3+ZfgnEohLWuEJI0/n282uUfiwLR
EjxAlzRHsWI/iW6mmAKxQtdKEilrRPrk1Psxw4bSV0e1sAxYnMxdJupIXIYic99f
qTFUNdK0xpHCvvDMbRCpMY5mIV3PGGGW/kZMqR821pYTr8yXckOMtAT8Vkf2JB0v
oicSzyD1/A3fwhah0k+Z+Uu/o2FdUzdUwl+3bp9fP4VK7rjtQfOF0GnzHO8Tyd4c
CVRMs2jvGZ+6cKoURcmhk1NotPSrGsjtRh7b8BAIowuIoTlAMZ8lqIpxVAbNSqm9
R4vznoXU2Wt4rwjdNV4S2e3h4bm2uEoJTwjP0+9b5YBOynW0T1nVB0ghGHWMasZe
cjQFPY6cVp2iaEHYQ/s9lFzqsZ6CikkCtDRZVQ4GgTIBuAIKgTtN5QD3THDf0i3M
Ev/LdsjO+LnRpEGiT6/ZmlZG100Wl1+BOqs/RaqTXyLx/2AvTZn6++MIlMVZ6UZB
FqVWkJtDKIPTo2PXgyLh246ESv+57a3941drCMNzRLB21FxIyq16QSVSXJm4Lbha
+cjBZzeahR2RpDZQBiXhuQhq9QApqvCkXwTt1W/kO8ClQrG5Lsi0pet1CiZoPPp0
+ksb3Gx4efrUA1dk9QwgSFwLCZ+dTIepvaYyni6SD4kaZSf2iuRBJueV9ctSwwhp
rnPYdEP5HkUnoHQmB1MjTQkxAbgQ0BcrXbSVzmR3kx2vXYqGF0TpQnmbHyYypyqS
KyVAbtqH8fdZ2lEapPvYVe7/EenyjhNvr4B7quhrdMU+NjCn4zSaKeRcRp4Kl/EF
yNGTMDtDYMrCW5ZOvTSgHOzNUngxXQMiJkrW+SiTPotTQRcKkeiWchhP+tnbGvQ8
zxiAEbPnQZhEvlEpFq9vySVtssuL+Nsm0KMU+tBAfQ47kW/XpBfT6A9PmsSdPp8g
mkmOoM0xbqzm7+Z5kQmGyi7PvcLiDob4UFMPMeah60k02ckRWnl+kNUqSsMAkGeY
7oj1wRANEnvtn+PkgTu5K/TnevRNwuDgZp/24PzlRi9ANTJAxu4fTnG3qujz4KGO
Ex5ffBjZdLXOnZHs2xlFjY33fMSD38dHxM0c00vcZZgBDoNO5KHSFu3ch4bCM7B9
LGdOlvHWdBm1K/MNFsi8US20/dy+RSpmV6f1In/JnTPB1cBllkSXtPcWKlHg+KlY
yuRyqec6mMf5YblroMsqNhNaVkhyiodq8J+AlvdgodQDhoTfUXJfMrWYyySTsrkx
zBHzGRCFRJH91+VP/6IoBzcJ5LoB8eLxLc7J5Dr01dS88fREBWqx6o19yRHZS3bb
ZtGSAT/1pKYEDJv3NqZDUnQkIHaJ4OkLQvH/WZ2+tokweNE4KyrnaU6g77f2tIqp
Sw1Ln1VNo4j7oncvZMj/bNwxdsv/Rc/u/k7xu9+E8GLcjBE5eA4Vf5ZH/fOGlRSm
YxC/ziKa4TximlrpE+jYRY4k5xdMNzanb5GObjNp9f+fF64Ke7f91JKkkCbVOs1W
N2UEu6uY+KWOEGiuRqzZa1a7vS+1GYky4lXZeHL3lP073O/O+tiRpsSvSsf/Eo5T
sbMswVUHLSfDzYHbGLMVbm9ZYtrn1MpJrl+MDaAzpFZpF6QuUKFga3LirrgdFw8L
gJtVpIm2N3y7jQQpYk7yrqPj8aDB2AI+Mi/ohy18FX82d5syK9N6QNAyaOyoS4OH
YCLZvBEuwQ09u/lv0EJTObMH7tgB5rAtPM42LwCWy83Pa1hvuIRssva8oA3a+P5G
oneLcnN7YNxjbOLB66UGWlnTvE91QihYXYFngD5mfZgO7BnHX0CmFFj9HQKGmZyn
dQrrxEYWN7sGemcCJxpuPH1Osp+nMDjpS7+fvKJh+aFX4O5kYnX8xcgNjCnkc5Xo
OfT/eyIAWAuSlue9+oB1l2uB4JtN4kqpbxXRMgeTC488dAOLu9Go1sRVfUS+hdMg
E/Q7gwUothVavBJqpEdMtkHu0Wz7E5SOfemvk2/SEAgj0P0owHPkP9MvIuOPvh/C
38lAzkMxOv8p/dubL3hgvumKCSwJUPpnjEO4yu6/KmNoWqHoHFmYI3HreV4LyqxD
AygK4WVY76S6glb8Y5FXmt+UQY8zzVTERVoyfL69VN5Zz1azkzXoRBObLy086/dN
ERoX3TDAYCCoU8EThZr0WP4g7I6YSIgZE3ezkjZWLcp3c6TfSP6MnzqwocjZ/m0z
q2as/dS3dtkQ3COLmOwid7HGLJVMd/Pl0elZ5K5MDY8vUgqU2y0bIY2x2pkSaE76
M3zpvO9wGiA4S0/JcRkJhkFF8dORyUOknPHMFB9Knnm9KPp/0qNngTkPQlUnDVA8
d7Mk3Xt5Om2oLyFOnk8NvmpFWqJHTXPqa1gaYly1/QKU5bkctzTBKX/XlnN0X1kL
p8RXntQQq/GW/GvnxroAzL66W8QIF9jDuC5Qq5YwiohZt+jWss3sd4/H3MOg7s48
iw54Yjs23licHYm0YLIZmDUFn9Red7H2Ipw8UweclJ3ZxxQwyRllGxSNWjmZO2J9
kktnfMqQerpZubXSSTStbo2STxulASiVvLS0hum+b8gRdbnIoDVTDHFGg80+fGGf
SL+xlaQUmFp+eV1HO4MMWWg3KaNVdBP+K4S1X8J9WgY8ynoMqSrgRzn+pr84pqYM
EUrg+TCnKe/nOZ6oWbvzt/LRNI93T8EseiKoOssqJd1/qt3oJaLI2xvPTkunWr+b
xHneWaBn/oRS/4x3t4Sg3rGBKdLoP9X9to0fYfnTfK3mDAjEbJJPvRW0S9EiZ4rT
J9dOREeDcrI8MXc5bHDWWeBzs9DwDTaIlg8zc5jgufX8YJDDiEplIg1y5oCqU1ZZ
yB2bhb51Xf/iFOT/zvWGccxiGB4MM6MNtrn0/ysPHUQgd6j0JuIhaB0oMEjTDjKQ
X1sIluWRbtZykhWWjC37ILA/llZjbPX3Str01U46fayj3p7342TMs0j84P5Pb13m
jH9M1C4ybZe1OyLrs+8f/1loUt1//tA3DiVBPJEjUhNZJRVAENDOAvNtgOctgO53
dqb/11pnYvAn+4JaW2Zd2+HZlO4orfhXgPdI3tVAQb3+6O41SXHkIGk9jMxcUghN
J5qTCYkxTfy5n+38l5ruaZsfJU9yheH3lJtroEcy/jkHjmkOFJHlG5xN0fo48f4l
386uflgvbk8s+o3GtBiqz3S3nW3jKuagSOcw2xgxJT0iuziBHd+gZv7PewwsI8IQ
ROq8sozIshMMgq4CJJRgeGh+P/rTtQbiCpch2XyR67n+vrYNQ8A5i3TmgQMW3nij
nVolauN2BYE5p80XkkBXbTbJo/8j+lcnJKn8u0CVx2//lWNw+Cet0lvZ8ydN4CAM
JCXw8XaksWU8uRhDHiKHlHoF9F9H/LF+UTdlJgUgeQE53D19qygoBZp2zveeAEJ6
nKJ65wdWSatv3HbUkINoDMM/M8zGNrhZm28jtvabyOeCcVDeyZf/YG4XXfPM3C58
sRSXweubYsCxktkC1vdJDQAxyRZMkeE2oW7IhKeJsCZ1B87bqQ4bZvlCCy/+h1Vu
j3ozEezvLpCkJrq/qVk2Uc5raD51mmAwVBKPrBcOaaVhlGk1T9ughVC6EubVdF2r
neKaXPGtqp7SnctaFZTioRLYlLLnobnRqgd0OXUtFhq2ejgZqiN9rpKNtdatY4lD
cJLS8sNoK1gnMzyWuhB3IbaU290XzPnOI9G00ud9yiQESrl49+Y1UfWJqizY/LJq
AxwCeNHX4YuVcjpkP9UqxJUGt+SzVTfhH3K3aWTyMdEVPifNMIduuF9Ehq0Y/42C
alh16Bf4qTzVYkRItxZYyaYGXQl/uY9nDTy3uJOQ/A2p1cNbV3AEb0/i7E3sOJGA
r0VWxaLh3rCIbEnceQdRs4/bKF/cHkzKpck5Y4wMeGpg1IyEnhTMxwHl66X9LAtB
+Y+FVrAPjOlhLq2scZr/3TTlnwW8EbZHZXpiq7gYLvihvGEruVMm0VKCMHWSXnRG
hZg50i96GG1lzq5XrsmcYOA726Q1rLl6NzzYbT/mrMF77lRbRdonwhsakEWHzePf
UMRjBqurNYqqSFTJviE0mPtU3gzmal0u45RqXq3QqsE=
`pragma protect end_protected
