module test_top ();
	nios_base_tb tb();
	test_program testcase();
endmodule

