// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B+GpqHOlg7NksZaWktpbVhU0ASjPEICkRIurGySOHSJuQdGdxpJl6wUCG8Hjm3OX
F3pdYFhNSsM6cZh5WesnfwSdgyyinJ5agOI5rkz7GlMWeVQhjL2dNWemvfpSXnry
j8eJ+8zFElr4xcSZZRlkgHe8TII8EPQH95TmEhBDLtM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2592)
hBx2gKVsA6IrUT+r7KuEtiT+pe1Jvk1AkHW4ekab2t5hzQ6mWKOnoUmy5Lag12SL
qbx/nMnN0OOCfdh2pcUK8bmRgDKsqaOjP47Wl4C1XK8a/M93YfPCNTXoKdOhcXMI
OFwZY5CLQ+a8lZqeuPegZi0azPnvHCV1UFAeVmUJFAMcRCQIzELzpx4faLejRaU4
Y5V2loSjii5iHUUszFNxwLgWyLVx1zqqFLUg//WnJh+pTNaUfFH+8aSqDHT3HvO4
Q3PIr1DseuPCe30j/iWiDhjdiDCuxuhOIui2gXIM5DgftcKy91ND5tuVJbbJCdJH
SXyt/BnTj7Bnrimj9Tf/f6EEzRX+IUUhi556WUilriZNrzSXREVg6BhqoA88Acfa
AV3nPxER8/l5w3wi5XInztS95vCB1KmUHlCXyPJ3waagpFtgUelGyH3E8UwUowqM
qNfwiSC2Z1GOocyJlK1WrB75tfb4jOMfTOaXYrzy9YlC8CdJyShg9ceQf2la27Bq
cFtbK6LTmqOJ5xNoB8j2WPmpX3r+di6ya84ErGRJO/aUCzRD7ILcxJVkqoNbDQnK
Zb4Q2IxUBmUou2nkirhLrnBk4ZN5I/wwJX9XKsXBg2s1SjJ1/jlS8mGKIPwtJJFW
3mPPCOOumtCRwiCtIT2SVdMpWr2KViBNL39RO93fAJ/FamBuJBfpydAY245Fz6//
v3L+Vo5ASV4H3FdvQqTLrP9GnWzo4mVCGCKQh/AVtAOQx8+LPte0hev+ZWhFnBUY
5//gYL42LQSIs64MbQnTMJa8z/UjF2peO7vfee+T1Laub9rYoUu8Bj2jxgDiCI8k
CWH6hC/42OWpmGVKc/8OJyn1ScE01SvvPS2qYr1BGXmWB2g7Rn9nN6k6wcEPyVqS
hflqbVjSVzsHvyyaTOF60e0sK3pH64m1AwLSnioUECl7G5tpfnO+aONWkzr89D3+
6UffYUBjzYEx10tXYTEnrwoTKJp5gQkGkfig7/c5z/p+vicIofS6ziYlyohpJxtK
zcbQbMDVyXp0fTna6qvCPf7bi3nEfFMHJMG3cZ+e65o+aIln437Lx+ILz4KNyYur
1tQ9mxpvfJ4sj56eKA9OGWRRbjY2wdTXIRMrplh2H0EC9ZimUkEikRvQ1g5wgNa5
0DKamErtCXOoS/KJ+1eVHf827XFCqZexNlxPGFBkoyG2vq68Y6uokttT1E0M7bRi
MbIEUj71TLq7aVgQFHh9ixbM/CVMhq1g4p7KPUIYD/T7kVJwLL9TP0sLVxOEovTq
wVlnLwkt9wNYqb3NWY26lM/m1mc5AvG8kXLRA+ZKCPHrRcWLYUW/1Qz+IeLhhir9
01kSGQlTiW2gQ5/oRajbvXszUhZaurwuPXzRS+0EM2O5vjkRrHV1GBO1+r1vduZX
V+lCZNpOUAnt8DI0/IB+NPhyd9r9cTmceYhIas38x1jjKOFW7dvBLhOjV6s5Jqlw
JtPEaRRwa9560JJVb3Ixm6hKOl8jVxCCXZg4U8BH+HLEsctLmpzBn18vayg95Jrj
9sHSMMwCcn5pGqSaks7ZAmRD4FZwJXzOi/ZuViOodZ+fINqXmq7fK69qWgb64jL/
t2JCws3Jvz712GLStvMGCOayd9iUfuB8OR1kj+RE9DUsfa+bIlRGJ5IhrYVANR8Q
96Td9HiOf8v0Ot5h9tHDXv5ECdBIIDB5gIYr1N/t22EVboh06dSdN7IJhAWcQJcH
eOoZ7v6WdjRufm2usBgkqYh79f4eyYMxvU3z34Yh7Z8ikJoglYjYXHd2fVStS/Zy
T7s7ziLaSt1KMDNDDpnLtYPaxog1XSEoho2Kxt2eH0lCestrKmg1uocm0GrXkNVK
O3nVKDTGBwqGAzb4qaYYk6TsVr/+yTuLUsRsv70qbeiGAOfz6J4qpaUCw0yLe8Iw
kCyaTrMX9UmZj+VDPqfdkhesosJMzMt2aKvA1T5EYyxpo5Y6Rxs8Ffu21hkig9ZF
+HK+wKOGTA5S5UHWPRCcTavBSTP0GrhvqtFEKIABRsR0c74yYGl1grLBbCdb3OKK
Sv+iJDIzC8Ed5Tc7xAXNXqzOyc258RHDWeVCMKjUaLHuYnXKsYM5AuhUlX+vJny7
cEAVxea6kKyqjUwrG66NBtLdnHViSLIA6UvYhCy5liIHhv47ZJXPYrjKyM53Oh63
QIy4t+6ED2O62Jv4W+FC5uouQTcM+ooKh+63iHd1UqjHQybHz4fzc9ZZj2E5bpC2
WzYYITeE2MKh1nPGGrpmtDr/4pJAGY+rNFsz3ZgHlAutM0XelBqaMsrbjNxe0pRz
COmM+EGwpp5PF8v29GhGOmq6/Jnw2wp6JNYjTG1Xg5dNNu5tlZYX3fCv12bRYsq2
I9k2TtA+hUMS0xdICNwFGX8Op9DiyVsHpJ9vkdpVe4a1fXLN1hyPh1luOF/WxWcb
ILcNicZ66Ge8o1dyaj8yFk8fCmWTTcYFqI01EJvzBJWDxBgg4BZLLmCx/rgVmwwc
967Pa2lksr8zc/C57qh+9Uq9PU/SzX5PqF/NhtWKKwNSO5JTlgK6PdxSUnjRoygG
BDzjTI2VckC0e1lWm00zLChZ9VgX6IQifaDQEHbDsbQK66/uuqZc6QqY6cBhZ15M
vD7vz3IoUS5THK1j7lRitd/NUClBxQHyPW8N7IoixAF5pDgVc/6Jcbnoa7Pp5DLa
S4Pcu4KYmS1zhToJgYCIxP1UC7lpCt8Xfu50wiWmkOKGqyxHhC/jNkSvwtc26piw
A2zJ0lx9FmZenmzldp2z3ooren22L9fDoHBedr70gBrZuqemhSVYI0foTEerXwKN
5TN17P0Xc+9nXTnrs/20H2RnY9GgtuGi8Ap+bMK+YsfzASQhaJ+jseIoXK0vdwy6
RH3FPWsfB/bSIK/s4Afu3n98T93CO1Xsv26y+lSRCqa+vXlZBeF2EPBB/slqZ7Lj
G9k7OhB5UML/FXcurweH6IKcCVmrHGeCyhU5mfNAwKU9jRzIcZoXrF/dyHU4E1Nb
auc1VkcqzPvu/vAWyKxSvpl06i6IUL1kWCLHPFQP3a0Oo6hHqlX980GjExTSd6+E
Vn87D9M2VjSsi0NFaei9nAy0L/KKWIFf7ymHe6N4tjMGLQOUKedeTU8hfrclaYBa
GKWu5UD/EYcOnAf73zxLROxUDXjjSanlPW9WXAUlDKqzON5xIe0IePz+ywU/D7//
YUW7OoEc3FFbOJ5tvh7n4bfmXved7u05kKADFo1d+TtTtBVty/R7GmHxJGBO7CH3
EpqG3uhj7ae7vHSDRCRfZhr9SJcis8oGTPVNq8n1zlRkAEHr10RrN/5WVOezza8u
KJBPoRjCMq1tlS7w20WpFkek5t1uefiH+++fn504xi54R9Oh4cvdh+CmhU737YpT
6138g5pw1laQJobHqWSkIUo5dLoHiWAQf19N6wB99fQxRuCno0q/UwloD4rMVS13
`pragma protect end_protected
