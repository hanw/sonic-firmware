��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z��^���X�C�W"'yt&�E<�R�u�^N�Ji5�^�,��������#`ڑÚ}#Ҟ_4{�)�m�Ґ"�J\�sQ�.�9[G^��2a4�SD�`:������m�i�	��2���c�?�Z���x��5�'�Dw�w��������l:���t�UQ5E]�\�{�&��U��D�4��
9�hY6�v��s� �D}�li��e�g=[f�bw�W����5xӎ:-��{s/u���e�W
�HAN��G�"��)(�i�)�=1��0�v����>�X�!�\=:=�kh���6��{�휽��O�e߀��,4�xj����>��ҽ2,��K���@_����GGq"?��7���T����;�Ĭc��+��s��!D����G0\�p�7�կ͗1=@n ��?UX�^��1����	߰�,S�}�q��3\���L�/�Ҹ]I_�������=ҢEơ�-�u����Ň�w>�%��H���b��鴬kl IM��=�lf����������������#�'���sU7��v���
��mۃ�O�i���J},<5��9�aB}zN?�H4D��v�J�]9�ΜX�lͨ�}d\�cܳ87�_�'��`���һ� (]M�i�T/��y��!3�_�R�w�W��4dj̧�?X�-�t�>׊� ���VG����;�g} L!-��ĘYI�z�z�IG\�V"�Cw<���}���կ�H�z�k{u�肹�ԭKnh��(]�(�G�X-Z� tW����Q�v^�������Ѥ�w�r��t��=\x���C4�	,]�9z;!I� ����zĚR����lVR�����_MK����]y���ӺQL�]VEax�L��ŗ�^M�He0IQ[�q���S�	Y9W
���x���(L�a>��uh?F�{�l��c
�(E����:Km��W��݀ȕ<9\6��c<<NV��>.7�K���b	�/����^�ʜ�6�J��+��<
��g��7BqW���9̙�"�_�D�	�f�:0D�9ޚ�(�G#}6�� @`�������w@j|��I�@?����]\�'a[,�Y��$T`��lo�.��F��vW�(�K�Q���f{�L�y��g�ų�-��;�j
�I���䰑b�R`k����a�`4c"pD����@|K���{�m�n�nMcB�U��`ћ�0���d�F�%� �� $bPR���&߸����#$"%Sh�� G1o�9�h�	����l�dTdbpr�1�a'�J�5��w�&��m�s�)�UnNJ���g��5J(�'��͢��a*��J�6W���N�#�G���d��2X"���LG5�T|��+�KԹ�J=Mh �2�����}��s#N�2|�z�*6��������*�U.k�p�o],����ʋ��=v�U��|&ʂ�l��u��d��ܻl��*��\����
��|	�Q��Ս�F�v��ɼ^�9��UXv�|��ٰT׵��;ol|�"��L>X�2yQ�C���T�k���	�Ќm2(�۪4P��p�-+
Dn�+����PD��䬨Zc8�J�#ǻ �Y,��"�at��ع����<�k%	S���Ѽ;�V��҉(����ϛ���"�٘�
��"��#լ�}�uoM���a�����#C�{���r��ƥ��)� 3�;��#�:xh4* ��@yb��0�-�b���ּ�<2�;3h���OS���Ǘ�?/{�ƻ�;�`UB�!���|��#v�R�o�5JES!�����R�)��UzɌI7r:-PL�r`~p���.���w�ە!�ގ�1�h�"/�i�i�B����-��v{Ao�P���n�q��럴��I@�8��v�U�F܇1��eb����MEyC�>;���4�cXr����c�K���L�6��ص����.�ؾB�A�)�SK�'�I�����5��oQ�P
���$��cU��C��]cA��L!b99Q���;�\3�-�ЀM�V���Rb�OS�������4%ï��@�T��#|�p��Q�q����3<M�����\�'�F�Q�.��y�K�t\�N�}O4e�F<;y�9 �h���	��=�s�&Й����E)+k��=
�S+/�?Eoe����eJ;=Y�n��%�'����,��M�=���ϓt�Z4q��[vW�0#5�}Œ�'2��E#�Y�0�ƪ��G2�s:��!��G��f|�VpSћ�wM6��^tK�zNzS��͇5��UӼZ5��1��GO�6h�M^閸*$k)Q�?��z�K���{�/��=|hK*�A��p��˛0��}�TLYkW��/����V��V�j���
p��n��j!>)h��b�0'5P���*|%,�D��p|�����A��t�K���dAh�j�}ܯJ�k������ܤ�|���9k(Z8j��'�M�Q�lv�D��d�O�w)l:#w׈��uO�H�ë́Eb#/0֤ZA���}*��*����78����naTu�����Yž�VT�������4����{@j���F9� p�m������t/�{g��։Q��?ۭ�N�Qk.io�7q�&O�����v��rB��X�|�2����<CF�K�Ť�-�dWEZ�f`G ����>����`���[�?�;?la��z�ܖ2�������xA�n��LD�_���`^&�W�" �� >��-�2��gC������ W�ֹ�iZ�WJ����[�S4�ԋf�}[���_-g�������6Y������}�O×�\�E{���z�gh��s��B�6��4lܼ�1���B��]��#I�'	�@b��ݶ��3ӣ�����Ρ�)*'�m���8�Gv�XC9\����9_���]��u���Kf�:I8���ؗ��sz��8��c�oLz��4'C��V{��/Ɗ�ū���Z� �n���(/�؁&+�h��N���@�'�<��3�2�d��%���k�p���