��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���/���K}W��v�!��~V �qc�H_\�O<*F�v�����/$*oȓ��qMr������5���jy;��.Xޫ�Ѿ�=��'S'"R&�'g�#�ʹ�]�`̅a	�>D@��� g�4r�#�F�#DC�{��p�i��y�Q
d�0�������mF��r��8�~g�����g�)"�ro?�j}yX[���r�����rRy�
��Ԁ�-�C��X�!F�걉-Ti���ڄb��*��ۼa&P൘âL���͏qG��f�bvE:�
)��( �����9�F4�$[�x�gJ��?��*�Zi���s:��Я��!�Z��J:���t1�eyZr�%�$"�����W5�#B}+��ݜ7�����mN�v����� �^x�MV6ۭ��+�u�-7�ɓ]���q>�aS�۾�/�1�R���k���E�1�A>�%|�� �w5�8���D\հ�-�/~����:���g[��c��E�SN�Z���_M�;�lEILw��޸�Ԑպ*3u�m�n_a�ż�V+���(���]�X��lZT\o�C�8]��~�SW�y5_�U�B�-����A	�)��%
ݢ��Ȳ2w��Fk\@^��X�?�Ðs�{��)���"j�T�D��pp�������$�I�Kl7�Xn����`�r�Kk�J���.�;� h�#)A�]�h�.�"�?�g��]#��K�f�/`6.�#	v.Gw̐���*_��JԂА��1�f} Z�MNj.�B����N:�j[\��8�&u�0}�:��<�>�MŉI_�5D�k�.6�M�~�e�\���T��\ <Kf��<���t����~`�&�Y�ҭ�%����)]6Y���Y�}0��(��1��4"�TG���}��ܮ��ۄ��dbP��+a����c�'R��q�$j}�T�㗠�gqi�>,>����+!$���E����b�)�4�:LV�0�T�i �v2v"��nti��3�mT��W�e>g�xJCq�-����G݆>xf�&�X�����Գc�#�Vf�%�.���Z8���IV����x�L*�n�JA�����&������L�� %R�uƳ��b�R��dro���n0k�S09�`��L�EpM�垕-Z?���5y"~���$�G��(}:9�A��S���i�[��h�2�����?g��V� ��̿�g+�������W��H�km//�z?+.V^g����	��:%Q&QȪ��b�]��^f`�h�
c���>�H7�
�?ޭb�3̽�8i�,��0!\`�ک�kJ)6���,�D��$\���c|�]6�y+x�����T!��A��n�$ǹ_��Fu�h��sE��}��D�s��	+O�V;���r,_`2�z�~h��m�8��5�z����iY`��~�� �:+�:&b��t~I�R.�ʪ@�¼6�+e�xS�F�@4X���t�N�-[�[��7�ӷD�w�A��	�ŰiS�+�:�ԸNóo�zT�Į G�Q�C5�p3��!��:��Rɕ�͏;C��G�h�\~^�����_��N�C%@Z	�:� 3�l�����qO�ΙQ�^X��e�A�:�(?��.�Un�?­�C�ϝ~�I!%.� ��GW�H��Q<6�������I@��/ȄtF^��^#�X�ғ��dc*^�4G�5tN+�Ǣv^�+��q|�KV�LLm6�����ñ�Pˢ2��=S3���Qm�-�6�6E�pi����F����s��dL��Ep�W.���,!��%����dm���2oU´w�~d�<w���młAKԈ8-����X���?0D��=��Ũ�_��oW��	�k{�ԝCMTۿڗ�?ʰ�&Y���b�۟ �h�.H��KիZ<����~9�N�Db�����a� �uցqr��6��P7*I�u��ů���<�o3E^ ��}S�!��d�����o����6o�f���2:Q������ƐTɞ�Dy+��\��Mb�[�r(��@I��v��r}c�-��p��nf����
��^pF��>�$fJb�Q�ŧ�!�G�Iс�NE?�P�N���Y���*T�Z�ŷ�;������f���j70n�����+}�q�h��4cFCo�mD���҂���>;<'�����!�D�xQ�ڤyi�!�3z<��)�O�����_7tA����a{9Rج^� fz�c�u{&�U���8���$/+��/�/�c@?+�N Y��]W�
ݍ�����x��j�kpˌ��P�ٶ��!6�" 1�?+�P+�H<�6�?j�9n�U`�D��<Q�(����;�4Jǩp��k�F�R"�������y
e�� 㫡���4��	'�ŭ�������(��O޿�6�e0�5��D��߭��jP�~�9Z�V]�IM��ѥ�Q��=�p^><��n��rWʯ!}-��͓6�l|����]�����a
\�21�%��~�逡�;�]]sn��/,�U�z������NV=���Z��l��T��w
��c�Y[��Fs�=)��F�v���H�D�����gv��tz@�\a����0��g
rl�O\�'���KD|�����T��쭸K��t�륆K��7�n��Ƈ����3$F��zVD,�"�Wr/X�a����N(7ek�b�BvTz)M�ۀ�k�d�D:z����D;�"Q˨(�oG@�Θ��������H(��~������3���Sz6o�Lc`8��#�x0��iqRp��A�sـd>��k�I!ePd�'�]w� "�\KA�q%KxQ�[0>�s`W�M�H�t����L���Ӹ�%�-ȹ�4�4ɘ7�Em��5բ�|ʸgOLw���E�������F���(�u�%&C4�p-Ke��"
����c��ߗss��&�P��R�|�\��"i�_!�4}������ٖ()�	��[���i���q�c���kp^�2g#YrOZ*�?0n�#\����B*�8؀�JK)uC�����*ɐDD�Q~��Z��'ql�8YŰ�F�Va*Ks����V�{�U[��D5�D�$�9)��۰�TV*2aђ{`k��eћH2}�g6ؠ�1��C��������FFC���ʍ�ڟ�2S�Wj_&h�*��Yn��[�RF��fg����g�υ�*2����c��)����Z�8���Mh�c+���/J�Od�My�=�f�	�
m�I݅��]�U
��z�C�5�'�����A���c~Xui؉���*�;�z��:O%��;f/ڮ�@��d��J~�aG���g�af-�W�zߠ�Fؔ�1�?�1�20�2aL��얺���DR�G�"������SSY��@�:uR�v�M6�'u���z�N��G��l�(o((��z�����6<<�Z��ɇqdս�������.{�B8���i�ۄAn��q�����	`Y}����Q���^<�n
M���2 �t�9��Yk5a>P<�u���r�霥��܎?��f`��?��&BS��eL�?%üj>Q �*�k��69�؎�%��z�<�q�	[��e�B��T �2��.�J{��^�G�st��T�;�
Eñ:e�~�9uV�K蛸�0nwr,A��w�w J.�|sLƫ]�a�6d�oY���b���
�¦��&(��Y�x#Sm�P�b�1�����R#yr����������P�Sb�����	<9 ]����̂������Mtǂ�0�殘ޭ%٫[,z,ehF4?��̈�@VQ4ף�Ĝ4	�"*3ed��Tb��%�>�퉏:B�q�Y�ݴ��>�� *�jŖe�o���o�D�B͠}+s�&F#5����5�W2������w��Bݭ��7}ę�'�0�2�BH�}̗C��}�w�`uj��$Ĳ��; �7v��t��G�{��ɗm˾��*eѷWQar��Rn����N�s,��m;H
�Iڱj��(��DU��T�|I2����r�th��o��dܱr@$��%��i ,�hQa��i��֩��������;��}�`l�b6������p����Β@v��% 4^�X �T�-Ȧ����l#ktW,M
&	�=1�2��|�$?R�1i���с����S"o�\�3z�WG��ꠔ���/��Y\����^H�%����P�i�٧J��|8�`4w�>����{.�dƍ9��?�I���5�+��H/)<E���%E�J���I�80�|��i�{9��pB�����9�j(�j�gg�?�����~��A�3��1�G��\Dԣ2���&["Ѻ�b��C\��Cb�ྏ��*��D����H^�@����(*���>
�'��&!�1p�j2���?1P�0%�T��^%L!�顤�#�ł�M�� iw��#�%h�����7b!յ�h�'"����Ou~����on9����~�����D������` ��\��
/l����x<�<�X�vQ��YG�R�6U\�!(�#2hԥ���8^��;x�A�=iD��ŷ�
-��\ivC7��6oJxf�ҋ��0ÕI�v���;Mx��jT�U��=����˹t-�*��r�a��L��y�9���f���em
�AȨ=�S�D�V\�����<O٩&�Ǉ�ߕi�C@g���rX8���_c�Z, P��/����Sm�w+�.�R��Y:]�a��Z �_�MaR.�s�݆
5J�F0�h,�s"0�NT���8d�H������?66�FB��}�v*��e�"2Lk}oL��:�i
*�Jҩb��ի�4�_=��
�#b�?3��#��'�P'`f�7�a�`��rrc�>Lpo��=0)(�uV%A~#�$U镾 �|�+���<}4���~ �+�]Ш�ҳ���'ttT���Ќ�����
PG׾۫�aW�oG�8^��N�c	5�<�<Y}������.{���T�u �V')�G��܌�}N��bA�P�˷�P��D�4�ܰF�#)���K�ap����q�2I���t�x&\/Z|'��沞����x�ztq2���u~��YS��cY�"�y�L��$�/�ٴ0!D�E�����B)^{#���A��=J�4��贷g��X�YjA��Q�V"�1�¿�}�F�G��������:u�ʾ�}oZx� UwG���͗_� �!
7���I�)��N�u�$ߘ _P�}8��S�r�b��3��0�́��n�D涴b��n���2�	�'���2�<k��� ]�F�`�Y����?��tႏ�)m��9�c��J��w��19�����@��ġ�h��3j��Ar��lk��FRG��fqwİ�e��	�j�rE�Z
�6
dSkAy�nGK�"�-QV�vq���O����@�V���|����}�����F�BI�Ӝ�6k8Ŝ�0��[Թ$����i�'�/��A?��G� �]�HS�P�QH��6=q����}�m�ZI f�so�~����>��{]����5�`�jܸws0� G<�