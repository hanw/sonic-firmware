module sim_top();
    sonic_blocksync_sim_tb tb();
    test_program pgm();
endmodule
