// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QavsL8/N2uhCFZz8Z4GxXHV/gYAy5PyTedy3017K0DUq/pTGQ1GSs8nslaRygxbg
S9aRDTaluMinV83Ngk8+vbAGCRS5efuWsbq3cqI49ZHvdrBVwYI5Nk2FKTx31ekn
Wnim7KWsmU7QeoEH3tgLVeoCGg1la7wqzI+0sii+KWU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9088)
Hj3yjc6wnRw9IjTcSBmc4cpn0EyFRxp3IimSC8KEgAQEWvOzUROoy21uuk+a2CHm
k0m10WWlkpnccH5T0u4O5leuhJza/7h3jLml1rehSHacn8v2OZGl4wfYnkFawWKQ
ak2kLLv+HJGNtG15pRUEW4M3/UmBmugiurKkYFnQUyQaNPbFsTw8qikAGtHGpMHC
xdtWvVz/AXGucOMmraM+UowKkH8vS653aStGjCX1DjmNb4lyOTumE4mAnpfOQz4R
DLT5fjJ76NQ2y1gNRKflXDxdzq5uTuTV/z7XRgoLoQJ+RrgLqr7VY7KF9maEtR6F
/+1QhquJFn8wJBd9RdtyUiQwuerznCSlP5RlrmTXpOadTx+jipj6QMRVV5aS0Wjs
UzHPEgDBN8AQTvJm+QEVyB88AhZ7+5MeUrLQt2OiHowEiVg16RD6TqJ+VIRfMGAh
dSUufyaQnA4y/vIo9GBc5l0HhhlWC6DovdDgjeHqhncpvoJFihO3c1I3zrfuqgPu
Ci7ZZauguQEI1tyQ7SDiYNkE4R+mjFCXPFgVp2ngtTpGaJ7PQm3CmsWXybhga7q0
kcHXdePOt3d2DZLZN8g4iQADjSb3ErqFvCgmfvLetOMBvcTCj9hkhKgAPVK3x7Z+
c9mU8zyK/0yYGDcFXAgGmtCQYIgcYvbXSHeqAcMeDFSpRkh1FD50jhCOArfdfA/F
m1ZWSn0r5fJcPsjxbkFfKSxCTySCbEIOHeDyDuhIkPyH0y05QCcOlAy00lIRh1D9
3rn0V48fwxsKSz4ADfsH8/VeyNWJJVWIUo8ILmI6VB+SlciMDCUXiOHwRRWfit2X
yEbjFyyslDANEHoKxFcOMkZZGVGJabC3ZXdLXGBqTHdcTLP25nS1ogs7eYb3n5pv
Up2QS0YxyX0KCYNqUkN5U8hbYXmjdIEdEWmLS94kclXDst2lZNLisAzakcupJdaH
+Rzh126X63CMH00tfuZ8/WELQBniyfp/dEk4P8mDrD6wrOB/ffqI7Ndk+8chxZeT
MSZQby3H1Q7eY9KZgIDuNhUZ8yB8k/lbfUu5bGVHnPh+OH6gpxxM9BroiU80RXW8
0KK14XVaseSwDyYrScZjXmmZD+0JdtNVbWem6g0ijEUzbnyMlQRAaYnbSgAQveXF
UlYoRgdGkGe7npDxcEU3ARglAMqAWt/6JguBy3qDJtrWxSI31rWE3tUQgyr4y+6s
EJ49K8z3Vo7uKeDQWOGIUkYpqQuhkZVBkA2It0QFnhTw+n0Csrc1oMKX0CMW7YiP
6xV1/NsMAC7YDqb28Gu/UWhk90bX+fFjwjPosEhxuYmJmG98Em9I4oaZ4EtKupUA
EPax7757dgTCXDNKEOhWcMnJu+N24cdqiLOw4r1Ijs2/9lTIESLlpS6RAwFlhovD
fZFlhFci7u97Dy5+YER6rqCHqlpUEoch6Dmk5R9EASH05uffdqrC3fa04FkwluNe
vE2J7gxsNyjVudo+2KJgbXetLYjxlXxYo+0vIToHnR6trkqcVu+cLyvF5e7Qva85
G5/Eq66Ww1Y9W+ayIGzDgG5Qh8TqCHZng2tWS9J7FdmpYCULUkPfwHZVXkDRwBXs
4ZM9ZNXhBikfsIQbWkrYdIYeS4lEKd1d4667GLC+yEnKrKzfs+cxpmL24ah7BrOv
l3GesVj2rRtjp+NnUr1+pJQrw6ykqbkWVoHzuxPw5WNsWJcIFeoLO5UQr2zRhRkQ
fGLiSO1rxPIT91ipeOVT81ukq4MJck3/PM47VtRZGAmtTqdfFw8imi5fk1gROV7o
G4LM5YBI13o0AgqTeKVzeVANe9cqw/v5Q7t9/tetAPm1bSqJUvyMFnDvv4C2Hm2i
fFgaHHF338f2n7wDPIzB1fJ3AURPCUwBaUKoQUbiWpPK1PD/v4lELG65wQcT1g17
UioY5RgippUpj+FHlQQ3rkZIB+qNikh3HiFrXj+8UwNpSDJiLyIgm4lnJ4lY6mGl
lO2BTHcQucF9H1dsM1fiRG5+NAiCwI+MUyl5vwGd/ui3qhlXwQi8ffu0Q1H9B9cF
pB5zAd1muXnwYduEa8yesrshYl7UCp+CYsM5bB86g7DbDkEf/SGXU93QkRlA9MWq
NglO6Xw/cks2ukyoaWQHFp79oBhZVxca2ELvInQbBekJfHah4FPRECBpx9Erg5bO
jf5zplSt0na8w+jN4p71mwEHPfMnYjHI9CZLiVc4acj+xoyTIhRbQNsRQ7mvnYhG
RqTqixNfSJnj5tasFJCGgh480wPq9aZYcK/zvO//DyRx1pa+I6lxoR1l9agSjgoQ
Jhy4erqQnVD+ua1M9AeFjxOvT4BFnMx6HVFEKDdEL96xw3WgEB3HAxMGnUuWL/G9
h3K13C6JenqO/DHTxmQQe7tqVWhGsvpjT5egP/rAcpcZpAF+9xy1b9+PXSTeQHho
0sFEOLFUoT0gNgMce1xp080pjZZn0XJS5SK6lkHi4iaglhUrxiwHlMWHejtOtLE2
vbUGLViIuljUsnbJNkkF3Ksv1jivRhHUT/u8zudsB3MCg9nq1kOaB8qn8mnM0cYu
vDx2hKy7DnygTbHH2+XZ2uFPg0oM66zMloszoShyEOEZw82JV0gsfWXrf/l4gw9N
K//CJuMRJ+dTeyKN2X2KuZnakwsEmAcWChparnCTILjxsfXiAmdNCklH2nTYpG28
TzYLEncM+lzaW7N23sEBC5p0QV0SJ8iBcuUiJGhXvIv2zcEju3zvbbGhv8v0W+vo
FQHDMJQQcr+h06s/3xtKsBsFtcToghvj64wtNTbvTQSutFSMvduL7QyqGXx3n8qG
bkymIaZKLMgkpNeOvK8WHJcGIV9b8/wv9Hiv8Pyl/spyCPP828zNjoLvLAxP+o/R
iOioyt8uI8OYx9U3FRu4H44FTCxllbCWrpQXwGtu0ujZ3h6s1XYl72m7Lns5rIwG
V1+lSlXCXx7+w2/2dlLuofMtp9I5/Z5ByZ9KS3HBq1IZZex9AskGSxK1zB8IQpN3
LRXdZF7ktKM5jwKIPU/4fn75CgAgNle+OAm4Va06FBQOHiHMgsOnA01bVh0eI/p2
fQGeK9sRGQoAWAMshPigrMZq1tCZULxNBooj4llbJmSSsGBOt5nNEZ3rF8uAS83H
V4WK0mEpM05KJ33Pib6B9LvHrM/ieGlB5BB4Bu9TT5MdgMYZ8sCqWJCRelWevFO9
nIs5QdmTZptp8iS2zpSti7FIWQvAwhnoXj3kKrZ8f0f/g5ypVupIuh4LjjmaZb+E
GOHiLDZod3uPeTrqMPQrAfRzcOozkB6prDKptV3+Sahrklhz6jNnvW+eOqSmuvSt
8yzZzEousHTQ8DnPbpP4TPEgq1KZT48r/loZt3km6Ef+dyWnCFmrN+aotqNGgl8Z
NAGrMGXFNFQAA5iPXqxJwbG/4U9LkkACm7I33rTH+JttJVfr6H5JB2QwSmXC+tI0
Id6VqmnFi+ByJUznSD9j9YDlt53G0C13m2uf/QCj0OZGm58K+0O3/AVnTMtg38WD
vvrTRN9zdHOFHLLYe9dpve8BZON0MXRYDxND/Dkg1WYcujVfRF6Qnfs4KyLbsvUW
efNj/psBnayKvYHMsU+9jBSEZcPwD+Vy6d1aRjtistidSAo8Uf9U3fiKFUapllGE
4xqGZ/8uZ5+hXfVYjEeqabG+6FigTTkKDgkQB/ViCGWhRJ695bHR6vhgU85SNG9y
w3dMNUwdNvL5lC1TkPuqfH3xtXt8KEAI/+S+Bi2SaoivUlPlXiGsxexBS7dOGyIC
biKZCYA3bBIPYWH1uMPXN8k91RCwnZpqCndtsVRBxp2eGLKupqZ0VbzFDktZEMdZ
0ceC22k4jgrb2EOVoqVHlWbRTtGx6aWtUu5HWRAPquVGgNptTmGhW4KnhI1FQOuX
HbaHHbAvkfJdEiY6v8JUv9crOWG91wXsNyEOhGLJcJpz4dyUQkQjRp0vKp5cW3BX
aZ0xrPwE5Ixi/Jz9Gniq1D6Y6l8e1OGRluTWAhGN7mUtwKmB26EpF9bAQVw3vZiB
e57Rw48hf3PMaL4pb6Wn2WnrpIWJ1iwyAaGp3dgS1LmgORDRE6unrKNAsE7D8qGC
oAmNhF+XzkOemRxLhDEZxoVeHtyYvPer7i02ICnGLSRVOsRe8/Nf0dSZVLJze5Up
9hiejiyqIAYiQwQMmEKZ23VMd2gI+JudFuGDgSqbUyMfUlUfo8atOxN+Ag/1mhm5
ULqcAx2ORKT1jaJdZqLKdjMqoz/1aQPk0fbAoLREITpSqH5WiZM91TBHTlvs6jpx
aqVwbwaQqMcep/BvuEfL5XGSX5l9zkwonbptAHa9jpRCdAB2NqLQkLbrlabbjyfS
hK+Wpjv+RhxWLxs4RNyP0vXCtn4ES6hfzqOrzrFdTAgOaZeEG2NywY7aXB9/TGEY
kX88f0aml2N4Mt//vhx3fiey36Kg9ENO5zoVVaLQIhf5YBqV+ZnKbh2jyPLYv3Wf
5IaVd5Di6dSVa98vnS/JZxOsS2Y6iognYW6gl5ucgwTIt2QPXHvsV3Nozo/koMJz
kvyQDdDNzIc54I8Bs00NpgUSkOySsYUkzQUW9I2bFvmp79BUDaY+kJrXbWZ/+9b2
/+j18NPRPywr/GvfscH0pBwkieBIFhf9x1MtRc01Te+75Tok2n2Fx3J2/9l/iKaK
VUPKYTUOf85kdXBt+WpD4YZG+MEN7QFGmo16omeBdYjuU9Cgk6aaRcSROfwV0qRe
aiYnCoZaLgtY3DZn5DNGu4tbceiRo2QaE1zHFbns/2NMfvnYIXSjRNABpuqypIfC
c6325P3YxC8GXoQaADgOYJw3/8jyd24gsbbCDRsidpqtnD1z7DVh+k2olcZ8WpR8
m8WDRhpp6+85XEIXw/ong9SGj+IXf45nqi5rAODTDQAPCK/S2DKTZX4BOMsuVXWo
wVZFPAqY7UmmtNpNZpv7rAcYVvNXQrQYlcKKQo3ghwQ1G4UnVfylOFuRU3k2NWtA
qh+BfTwyLh56Y+8FTxe9yqlBMqQA/ntOibfNVgKVka90ksO6LO++iI3GysRxaJfb
G4dX9+0INwyYjBHjBXcIKliuqIHnpi5TK8zKG4nvEm+R2aZbOK6hS9QRWSN/4HKf
cOj/lBbew/1z9CtT8RUOBU7CXg8hE5FfXvdQypqEHa9nQTcDhKNdk5Eg0t4eHLBx
+CnVwvPsNOK5UWow3g2Wq6/YAaxLaZw6AsC7dmVPy3klOY0++KqvsxD23iIv/0FN
crZ4uUOPgyZddegoNvi3eNPnXSDe00PS1CTP1yT1at0Tb45Iy7z0MS70SKXxkBeK
Ixhngowf305KnIh2kNiQ/6z2cmNhiM7HA1YCAuwBLWTl77zqbJyhgthXCCQUD0Zf
YzLOH8c+M4N1pz4RmJetQqP+X7CQyUJPDvY/RnzAT0bxKAp1+a8GNdAVcae7sWly
20KYo8/EE/UMshtAttCcuhik42GSEhrvh8w7wNOl/wsLGN42BYZ/XG6r8I/hCksF
pe4FvjNdQ421wpMqYiRj/u0wfwacvTqX315QFi64FnhuUef9h3weHCOeR6uP/n+I
1TordE1ZvyoLKFhGqsrv1lP4RfWsZq8stp8QVDAooqRf1V4EcXeD7Pfs+pjbRhUC
pbqczp9D24nty+aCLW/lBaeV9Y/gZU3B+yKxcdd3Gf9FJmdRcC6JhASx7McTZur6
PSyu3sUgj5JzcQB+ypdSlpbarV7+IYg8A6gx+mVu5639vI/bdnmRHGG0ZI5FpYwf
LDPilb5dXtf6RT4LaGq3cKt94/x8ONMfBHYNdDf4nI+ztx6HhFhMFImS13I0E315
6xF43fBLG+2qB8+ixb4bUd/993g7b1CCiMvjOcFT7jGXqZ/fQUwWqNgRcWl7SCo4
kIUvU5OvayXlRQ/cGVv3st5xEKBZOaHXPZCuruWDOSiWFQnL3t87MfRDsYBaQdGX
fjt3T/g9oXjnksTrrnF1kRtAeZK4xqnT0TiAm4Xo2zEw33W2HzJ08jGUet/eHbr8
VNRvk+DV0/GVb+Z8k2JqITz2hzwqRGVGQPvf5UloOlKO4dwdCel6mQimqbi/WT91
KWoL+AbvXknIbJSWHWSAirFDO7oz+E5LNZNdlttLg29J0ru0Fneb5UzdvSiuOq8j
QGrBwXi6EHnQ3z1JUbT5h+OwIScT7pLdDVABBQMjCX9jAEA1qWb9+NVp7/cYzekJ
CtfKGlaJz5ZzWf2YR9m3II1IuByuQxQthd0AO1K16FoTAMm+Ntn2o3gR9gbxIeVB
oYr7g0udIgjLNQsG5Y+7g2vZzcpCm8UCg7FrU6HcYIdKq1Ggq0Q/IM2p/QBkGZQP
3euiS5fBZYVgzNstnOsG6psapeZWNMRyH3/YuLKqShhw/vKRU8Dh2BQw7/qo+F8W
biIhEJT1uCzWr9aIOqDvXcjC0sMhE5BFWlPMI6yS8nmHCSF5iiFo30Js3FwARERf
dlQ4CKiqlP+AVbQoXhemZcpskfyXfD5/QUPnUSW41BYr8UvN9TdwGSyEniszfo3r
tt6XcNpkkUVR2lC0qrUkkzJeIiTCsMRmbp2ymQ/1SBq8Nv6XkO9lSJCsOwhTGMLA
2Vn+aKZ8zzrq5c0A2+hXcbEG0V2M0s+axwgdrOJzZjbR7zS0ASzkcO7zpiHxHXEx
ZUb5R3ekNxVS5FGzU5mvL+hjWt3pZD7krMNG9P0wr9+6lkaRLbeHVdKoaXSsTQAf
5WrZT0V5YgxAMJtjTfcnCzPh74+yNdINrlIX6T5tUwtZ4GVgiY7iDWTIjVIhfhyz
FAjmJ8MaJDR/5sbeJUpsIXbcLn9EDftAmpqAMyXprc9FgjQjhyFZus/ZDHi5845R
GWBMnkgsRyV1iy/PBODZSwL+Um2zXPiMmtROwSIwifmvrovhQoq3tdXrE6CqkmFp
mJZRrYjZiIVbNwKjDb7LWwqzJZ1LFNCbet8frpZlEqLJykz5RgLR5P+NVjI2YBI+
J7z+wmso+AXYDr40AANSkXJ2j2uwlVrKJ53Py77FZHScDx8GQqm4bQBZYn3ze/7f
84jgWEMH5G2EhuOB/tkoNzzqbreU3f+Qf7IcpC/oaCG8ZR4q1nCl2nH6+ET5jXy7
zyIJLqgiEbBCKG/bnZCnFWNWm56ifzbqVMA4/XKS8LpWTL5XEo7cFUxJYbNdhvES
7tp3od3YL7qERccIRw+qCcD+JFzh6zzXdLKQA3Km846wYPZ/CIfrOZ8DYd/3NG5M
gBZHZjEOgGDJQNQ6DKiYw1XZTANbczN8AP/dGZVIJ9HlrylJq0L7QAXwIzWGbBJv
JesCAEP59cbi8U/epasd84RSAc4XI8gtA6/sakL9BafyOm0kPP1Fkb62SKNqKbl4
jxrJ/HNtE5YUlQgtbcnVHhWAJ5xZTXkrWiSKZ93DO0oxgWyZKucBqxCWR2QpB5nR
shOoK2uJoYhAXGNFoFYBl3BHrGSG/7SV8zVLwE4Z4zKclnCeS62ZQCVWhXLXEAF6
y0N2SK0d4Z9a/aILM3wucwVHfN6MRyaPFGEosNFAuZIv4A8goDnNTEgy7o1+nABz
0QTNHItq/n079RtNiHm6nSCC82SwDpG/5yMExzbeInfcxAtwxeT4L0RD6SjZ5YZG
DRTPhcbA6iEF9UoY+NVU9lTYc1hyTNvUQ/HnI0gU4AIGYNq7UCHm0vlG1VHWsKSc
s+Af7fxoC7WKCKt7He8iv9Uam5KqRV+gu8YEBJ7q6xfn7ZE4nRATdlGeKvx7Yxpr
JWS+DYvTXxcQ2ZUhTcwsBr0W7YxnK8Rmpd1rOXFZR0rNxx5KRP+2PSdFw+ctSjka
wD1qPqp6UDrGQ/Ar+SyJ3UZ9HBfQ8k5CCtnOQ7XL4TNGgsNctl23lF+fqhKg97kU
Ck9epTKSo4enO74IIF8QOX94Lp8N9QIwwK09S/8xAvVybpW8HeQ4iQaoHQztf1kd
RuCeMSb6TIeY9W6Jve3HOS/wMYDeqPELx2fDZFHD4mgMbpAo235vaTioUqzhNcRq
6EcU38WfTp/RORU/KduZlad8eO9ObTHeoI4kMSO7KBRoO8x20CROsaVwCvZfiIo1
wlythmxyRixS5/dCWGyQszalZ1A9ChUQ9+DS0gjyzWBZjOrHG4/HNegURzVWgaU/
4u1GHxKVgEFt9O+nbA7ZX0ozfFXYKzKGDpCUUiVmaXyHK7wuZxCxzQkyR/i8Je3P
kOzLGKFFmVLm4iX5k/i5GxOKl0v1PfiGs7XS9kfNizkW3tfWlciE2P1cb0y9eTLq
A3t921UaJltIIbDoL9eD38/22LZIf46q7Z7gM6cNIlksUCQH4FzLKZaAqSkYoknQ
wNwqiXEP17VZVd460oktL2yaBfZkf2vUXKP01SZ/54g0kXj9QovOoWPOby2vqJjp
KHoBunogsWPQdcYBwwd/No8aZ9UXPr34/lrzTF7F2ozIXJndPcmsERSlf0vnvgQd
zPc1eL2cg+kEhll0YbbRYWcDpiFOt3jbll7RuagCMdwkmnTWmRAxhtuMBaAVJ+/d
TrRrzZpFdnaUHyLyQpJUX79egJyzDgXtkLEsEQThwtTfamOcEu66Wz4OxApmjla8
00DJ8Dci+qhT1lSjfro5gdDrvb+PwqaRTLyl/MxsIlTReyRMc3FS4vgBZA9c147r
6qDsSQXs6lpeh+D+C/s3Cmon+UFYvvnMBQknYjAhE8BLJig2tpRl0+Z3CKpRsi6O
IqOWZr9tICUHUrDZD2ZuEIgwxIp/jfam3veWb3r4+rsvfdYOVutGO4bzmURGS8po
t422Zb/8NeCX0i1w7idWSP4vxiJiyJuqOf/s5DzpRXQqeEPFx+DpsZ4R46Abnoj3
b//4MYya/3IyoAFNR1aD3njV3xQFxIoVzYLfdGfnDBMcNIbBCS6JzTH40LcL1M2K
eiqGw6zVWa9xfyAUNzLlK2B0NrsL00EjUcTCSFHTZndBOeeUsCsGOuvM0K/7UCfE
PBxujdCDQhcVYjhJFNifQRPUtdJY6IB1cX17ElX7Z1ttJthfY7Ult9zoBDUghlG5
qhylh8UuFJbusvb9PygczGoHmnN/3P2ASLBFAY/zWMfR8zp8SRBlez/wRSPKYFac
zEt7SKcJoJjQwqRTok7YA62epWwkjsQu+iAL8VFpzL4SUPkT/Sz9zjO2DtLhE7zx
aWkXC178lCjREEKoEaLE/ouNB/B2gw0r7wWkyK5L88uY5PIJM3jlwTYasWwDYeeD
yK5KddGgtxxS6g1JusQBqBqkQtaydoepWtYZxI/1B2KnIMatFff5ntkBoDqkEr1u
eH7aF4C6vgm8woqut2AgrJ81QaYuBzDL8SfAbuIMXjYCrc1KzlW78huuQwztJnqy
EfEg+bLZPIUcQRNr96yrufAEKzQHR6pdoJNOwBuqcv/REf3kz4R4oLjqtu9LRj3i
fwW3h5xnP8k4yddzTAq4iM338JSpc4qCA1B5HHpyWoUMmPCSMy5AErX4K0+Ay/k9
mjB8a8MVSyH97ucUkIid0Zc2sBXvxrVw/Jd8JTHWdxEN86/pSrD4WkA6RWjK50v2
1Vsd9Nhc9SEPKIfkYzFAeuth08mauvzbm51zPKikJg/FUOC8EbFGGQqZnaZpEPpP
VVu/j9sZUwd0/E2pAJvCS7JTDkkPz6FL5l/aY6tuuQoO92qHeMFM3EH0a3Y90/ZW
Sg7PeSVOojXXjIERENhfwYh24LUN3BmZLy6xKuCEUgV1vcztgZDuHIfWYpeBxjM8
2MS9ICIKSjWXUCjaf40fDBqo+rTdNT8duhbBew0xm4nXta8SvM5b4dgeVJYomRwz
WXfu4iXyCYWnMDIG73b94ZJL53558wIWN8eu+5tAG0BC04JUscMMDoZjdzu/UaBM
AivQ6EXqEhMVGzkg3K6hRCzfC2pxuxa6pRkSBsH6H0bn9vTfuG8ys4ezVSL4vYh/
mEY1Lk5GL8sxBR9QjpxsMwgFZF7HUP7b0anjn5GX9NwO6lZnUTshmQ1HVL7wY1da
AVvK+G4YY+6PTZ3fIvIjY/D0lgtVOO5S0LL00BrSnkTPwtfjs5BK7jdJgWq3GU1L
XVWfcIKDSHQM2vdBAEkZBq4PtqhGpVTPuuHRSGI47bVi3WzbxSNMDJLoSpEk9eFi
4qhP7fPUGIj+QSuwjonqEoRXzzPa8nOY9lTmNhAc6dbqvzkWZcq0Q29aFjyqhbCS
Ay4Yb1JIugAQnmTegC25e6I1Z18/fwpu8rr0nZYG4eMlT4cMioldGrsVLR4GxKPb
NYggw1nJJYJjxCdVF22JP2RCNX0nkjOKMHGq0HgRlYml6G41Y6S+ZuFXPd4kPuyN
kfUm/wRQEfxuk3V1LEtjoK7OCLbAqVQtjUqPP7I9n1qNxDLZl4oZQDrTwwVYdVz/
gzilC3MFcdVzWvWMgzPnHkdOdgvZ5PtcQI9QR2De+kIy4V/9HdgrY+9QmuoYcmON
N8bMtk0Cf+WMYqnnh2p4wwdaDFGdUcbi+BS/0E5Pu6y3zl6gJyHXZgtiLO+M5/au
6fCwwiKDOXddUK+jD/ywG2Xkyuoa4EzMMgusIHMN2bltSuFas9xryYOSIaZd4Fm5
57CpE+oX3Yh3/Q1Zzqzd64DwyJiLmpIB08xT/xbrOnzuAkw5TKwadHQW9LnLCeVr
G38e8y5ojPTO4hLOD5MaDBt0KFCVtlofkV9l/XRAsZSFMbcsHBJOSAkreaU39ZqD
XCy7CnYI5dijQtkOOfVeX6W/K+q2rhS/you3CJ8NJ6QSgtpdBuhoSrEPSixgPU6r
WASZ54GVtwEWIlDImEke/F871yeKTigosAmk7aeCgSo+cHHaRKgx8aFaTAFsqmPA
SACFgkBTrrSPH6xUNDtDvAQh/kAvIoSGMDiyWxSRUGNC/qOhCDn8c4Hb1Rwamix0
6XgkI3FprhiPwWCoFJ9LcCtTLRRg8DAb4SbJsMSRiSYuo+K1zxSerrR3+LkaBaOz
CvqXed+Gw2+OJ35FuerIkdRk4suvQM9MD53mK62MYbcgLUyt5RYMlP+S7Xxhlged
hNqgK1MPf5dH1Qaz7bOhFG8o3pWe7x9lgV042p7BPOsAA0KOQhJ/Du6vM1WPldBg
A5Pjmd/eQe7h3qHWRpEDDM1ZzsGWXxQDZl9buLwmLL9seANaqTHXFsAd419bb4pv
hcjblcyVappiYuBtrx4lEyNve6dhFb5jiX9QuJw/pQN752nNVz54zA266A1Bgtdg
QC0KL9NSH9TvEDKvgtbUfIp4roIdJKn0xbtZDpaaykCeB3bCtot7fip3yuvzl8ex
wy3SUg/ot/NYK4a9eVwgFeSI3OJgxq1C4rYRiBZyu7M2kNjLRNoSiOLcYFajoeGr
foBz82Dqkz2MFGqaNYYzLL/nKdwOD80OP+wKiCISM9CY2avY/Yx742wrqQyn/mti
HWP/WrwwHmCDb3r60FR1BIiW57J3Qu5Rm1IFQrqa5EErhLjv7bmCNCa8pyzS1vgD
D3/34e35fz6vbEOficZ0F+N2gq3lKSb7NdoJOkhnnTVa/5Lxz7eo5rxrgrGSwbjR
hdWady4Q2esPdAaXuDpGfWJtn7MHDk+LfMLTrpGx27e95qiivM/Klos2qX/ZIhn9
qShHmGgRvztHHaf1p2YqjQK8s2a3v3/n5Rab0ub7Fq5LxCVfE7qzMhiHt0RMvZXn
9r1Kv5XoPTf/zZ8A1THIvpBGwvApuPoezDiEBoOL6ZdlikuVnPUZY3NtMSDD4K89
8wckzG3075mXuzbTCsITPZeibh1b7Ejd9Op6no83VpUM/blUMIsFiDhhzByFlv31
9weII9UXaFskAthCTh1PSghzar7u+9B+plh2j8OrJ8QW3CV4rvU1nCU3TwsffZbr
iQ1BUM5RPsXtehFqkIyBd1aLCGOH53LOMxSLPqYD9npN++91tDL5mHLqn5Ml3YZn
3AYpWQMPziDTqi3TOm0q1tAKEogbtzQ77seoQKodqacsEbjrIogWzLKlSaRje7JL
Nm3O/MtApOIabfcVtFPzaS5PPbEZrqZKAcnA5c9hLub6uhWLGf2pJ3KI7RyvNXTQ
zoM2YnZBfmqRIosODwwk3seCY4VzIeRY4hJp8J4V9LLfbN1jacuWFYU3nlY5bFet
9n8tuQ05GS2iKjqBot0/qA==
`pragma protect end_protected
