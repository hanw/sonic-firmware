// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NG5nZxxGarYrX3AjilBsxE+m1CV7CkWy4MhMYnLqCWJ+QsdPhlQDFqICPQjb++02
dW8FPUhFZktm7Omn1ZbqYLucO4+MlI2Hlwn6/CrWRHRWtg6R0MWupwarPOLDLjRH
TnxXhIQmMyIJS3tZoMz/pHonfa1wJ2HPwPF7ttXPgr0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11712)
XYH1UGMW0xwvzECa6pXkJd/7B2MeVys8vjZT95A9ufyoPBjPiuelsO2jG1o/TmKC
dhH2N2OZQlh0pmwfWZhk8s7M/VHE/sSYMg2+zGSXtxO4QJXVMCjN2eP2M0/ViPlk
YxacVuUxvtIF8yFXMFu8no4Co4ovbX+wljYgEARJGiQPjMwjgbWnH9prr5qeGLV4
UlzQfTPFb1mi4HYWf2fcCkca09TLtfD4YnJzTHRHDz+d2Vkc48wMd1RfofHcKQFU
540M6nqdlVMOwj4dhwTBBsuUj9IKxKeRXQkdqsxq7Dle1VyF1fKVu2Lukq4zz6P2
yKD6NFJax+kk5d34iJbbUYkstimkOOvAfDArxfmYuvnjfb2nOz26UAuAYyPG1nNR
id8S4T8oEEAfRNzNV9GNRYlrX0em4fraVmEZkrqmNYCQ2fIh14k8CU3YDVix1lr+
i3Mv3ao5ae7Hx10nWZl4kgAP5j+9rLTtGfn56SA9pkp+JwrbBoYBBL9yLobZe2yX
2cltyIiHreoPegh9vcAfB/nD9Cu8xpVGC/3FXtVxeJtvwEQRIW04kRJZbQUKTGH0
riT0Pr++6gYOYi7433NDQYej4Pv2LsdSRSUqELYyvEEE7YFTAEu5veLjTjQWU92K
/Sj4w/YaFSv1cL09LAwbGXKCaCUV7K89Kp6oT4wANi9QtX2B16mo6V5y/pLOCwje
Oj+BEQXmw982bFjalP7vkJygaOLDA5KczotIpRWN/Keix+JOw0SDYFm0Bg2ujE1o
q/UZGnPB40p1rc2/Nm2kF4zhuJBO2MFY6e/M6uHWiMCdGlTaRSkFfaB0Ugm/HXL7
Kxwc1wCIAAL1mHtXhollaj3BRqAcH8MbT7felb+Ld2hXAjzb8wkzdBguhuzM9Nwx
6SOgNtJf6eTdxPxJm2lRwdMhEcN9dElsl8tTL4pmP0KLh92eQIbphw7YGmYKUqaM
Q5a8GYtN7SuH7yM8tPyDv0pyBRbKCH8oCX3uRLfomw9D0tbJn+o1sGVKassDF3Ze
3+GnXTPQdm1vwOWBbh7Iwm0ALd4UnKqGQrxNcyjIO+3yr4lqYJmZdUgOWnMzq70L
Bsnm79gYNuwUUCWEqD68f0P21UHpsgIvXmFVjQ7WUsl/X+0RnweEKRCufkfwlnrA
+079thR0kspMGyCr+WolSsTzwjmHJIGGX/Th6RSq9dgmUZyiy2z68T5WgdiJsyTa
XtcuhM+QbSK+K55YiPi82cpVlg9FKkQevFbctDyXc/kmT4XaE61R4HaVX7yx2MYz
F6Thqt7QRHZBuvBnR4+nlljuA1whAsi4u7cgYo7Rd+mrS7KDILSeoPdtma1cXz97
ZcTMz5Rt5vJnSOvuX6+aF+J+lysTV1WuJt6gLAY0N3tkY7+zYFVDIl0dvVg4yU51
iBPXCiTMeTh8fsVopR7ctZhDhUiD3uNQzWVYJOerTswGOjFbKxsxQv5nZ85YUYwc
uhn4SO/8twNpWyUpHtfvWmh2e7KNEEAhTU3HHnHOJyTLN7h9fbR+gETuFzkjchZi
q3enYb3WIAAeohb0yD/Q9HlI+d7XEJhLKvqtOZyLlQ5u4Io/wQOB5mb6o5Qs65Fa
2AMpU9T4/1giLnKF8ICjeBSdBh12823ZbubqKl7d4g2zayIU19PRDRdq2oMQbHEy
3qrhJ3ehZvcyoi33mO0Xer5BsmgbGaN/JFH36vDZBRKheLIt92iOEMbAL/VtntaV
7azAW0cV5CLMMeUzFlGw9jwj8WK7ZPFa5inhv0TNVYPgtJ9g8CaYNdhmlLxM3FZ7
3L2u09GjpB3c74wEr76MtvV9FGgzjq7sfaTO1USFBYHe/fvE/pAgpNMXNDjhsp2I
rUVD7oNFD6Z5EoMwQ6eox+U5VNiBKqg4JVl34KCZcpKhQPdXaoQOWHh9ZQZz9FoY
Gr6as+wZ5U2uBilSCu0x5z4eKLkBD40u3EDOPuTIjOUqhqtgoXzuXi8hO9lF5Kqr
321JISoYJ+ZU1tylmB/fAvUhsA1NsN4AaiWjm3qAzDCa3SnlSyhyIxfIrP9bUJcA
cFmI11XadrXn5Ktcj28mDhN7vx5kNC7mu52Z33gspA59ir1q5YXXrdH/DyqJY3TB
vK8MKRABbScAJF4vy8Pdx6Z6TGK9Wq1PpbrUsFJHfTbg4SZ/j79hLfYo//DUbEsK
nWt9mlpF3dThHtLvJyCR0AwCHQ5LAhQE74aEn1bc9kkoaLoVtCNa5GR8rGQRBPDn
TgeHXN9uTM2GglY5RI58mP4y3tpLFVZBHwwKbbeZMEksiKpXUXkovWOiEBPJoVeF
/EwsNYxBk78GA0kStcipNcPutp7xdzHoW2/pJZJwSKZOLHwAHOg+cwbXUSWSlYxU
PeIFM6gHkBP4Te+EiXqGp4yMCoXZrJJPQaIatWle0Xe3gaTNpVwIxWq3sfDoo76I
fKMn3SqQ/RXY6RM1uuvNw79dgwXrledNb1cvV70spzUmlkP094U6eM+546SUehD0
97J1aWX4rUm+LZ74l1ikqeoDDc6QjqIFdKbvSSv0t9HTZuKbMXtePw30vvbNiPuh
28ncOSEuImJ4jBdV26MT42jdalXzlEj4ULNpWjnkh8MxLSTvlZSrbxIrRAvw8WEA
GitwTH+jeIU197tInxFmFOR+Tsz+oz5ghxKbD6twbrM67lBiFC1SXsAiuI5rhn2A
nH+n+QjiSXzUjy9mRAjdoSUv03I9OyZmlI0fnnC5HQX2BXjGwhgAWB9N92qglkB4
JKYdLRTAJw3+vrXJjZgKu3yV4tr2qLxWdJbefXFnuNLjcIfV0rc1ybRLefW7sG8y
pQVd/f//r6q6qJr9sprdQBjeudKPVVkySZI75m8fcw65H69ZXL+9fXTIZ5n0V+Lu
wDGW5BT92Aw5xq9SyzHTRXJYBmJShyiEY3EFT8AZYXAVju9MjsiPOMje+deyBq0G
B1eKIigaT/aSPxYdrOEhlXd4hx088+EleNu2lDjKuk472LzdpkBdEygzSLOwJfj9
SoyFU09aNDbhM1s0FuI76mK2AARzrjKF7cFy+hiGywHFumI+RDhj7DMcYdtsMgIH
dsdYnDK8YzfExIL36ILmrTm1dgVh2FrSp4P4AvS7lwLHsAMtHEU2EPcjDH0mV49B
/tdOJl297Qu8pHvIg5ajF47BXFnHC6IoNroP95RAV8xl3uVBlc99722/Wr/J4YO5
nopkVo0rcZYCD1LGjWeaGMC/2+DxHOtPMwCQQ896lUfoFbRcMn7m+ny9L7n2RA6U
yows4kjoznGb+9kujHVcqH0V82UEC2HqumO5HEdmqj/DTlS0IKK8cRExMeBaUZVi
BJ7OkJhGZLJgUBI4roO4E5Nr9rgOhMr4pj5LzNoua54ydruBFiR0//t5b7zTEbtF
l7+ce7552dw3WKcqClzNuAxBQB21MU5xBH07k0dZzl1HkQXDYWV3iwQXydQVeih4
DoegcEyFi+Rhpgtm9O8v+QgV0q1qfsFpnC2RvIrwMQbOUCVvxS8xxC+lJA3WZqUE
5aFuYlFkOvasZ2WMzrhRChdZKOefzJNjhEGa6k2mDnnhfgC1x1+r7JGvX2ZYbZvt
SAlC/QjiwunI0iYVh9yG7wWhgUI4p6XqS5PRL1wi8lxP8fE+RX0WZPIX562myla+
AjKMaSnBiNmO8jsKyARBocfIdqCr65u/Fxa7LWRBjNdGq4VAw8B124WLJOZdK1CZ
oF0+Asnf3+MUNhQ/ixh6E5XVATIMlnPxoJNpfuBW6zWzBq5+p3IBoMfbxDnaMyaq
SYJhjIRTVqtapNe7lwHAAY8lH1UjQoT0qNBFIp56ZoNBXyhV1JsUcPtQUGKzpYud
4G6itAp4eY2xKv3Fv8cSvKR680KBNToYhQQmg3UZ92GsTVrFUM77ojuRhS5MNWGb
b+h7DrNo7Wi6j+AKzUgAfK9WDxMFqA2MAgJ5zY6G2X3AUypzZdZdtOHTLIYWBcd9
QAwwWYA0bLEMJcfCLcQU+xmQ3kwQdDe5N1KWpSi+WRYvrSHZs2QPchdzdd014xWa
j7nZD/RbzDytdNfVDElXmril0ouflmP6BrLEmZRSOMW2u2EsK8GTrkJds9ChjtT7
F4h5OTnpWVd2Ivr8eEQ5AqW7jXffZcOcmg6QxgFlG8RQiOfCr6Uc24qathMPUJIP
6vF5sCgTVwB4G8Qy6W0jC1VvYa0KZ/rqC2GKkljCDaIlCfY0wIVYk9IDEb96M1wI
OJE4TSLCBjRifANjFcEdqZyhJLETIl3Dl4Ey7OZzAwV8xJ37NDVncsw38PRI+ksj
amS2QiVDao3dT5K1O0C3BR0ypfNd8zk+RSUn0umcjPxfytoFY9j3x723Yw6JSKr1
FeUYFAX2P6rL+/+SkkB8K1VgxY7J1fQMEyd4jgCDzu3GuO3VKS5mdmrV/sf2CuGR
QmA+KTYfiFjaKUUCnr3/su9/tmnGfcp+idfjZccLRK+GbkLsh6/iU7iMlBhZuKzZ
Z+OrJftWJQpnsaBqDbMyc5wnemIboTL8tk1vfjb70hH2uQvOaky64lDEAtqrUh0L
Jzz5RsNvo1p/yc0LawqEkUPMBdQvajHi+gWOXkr4VN+7OzkHq2F10N4p05MIUe35
nvrckYa4ClqUYgt1DA3ywAcRH4wvxm2XiXh1cLncOij+UE4mNX373oqDcHAXiuxA
mqHxTyZbC8KD2WLqsoYinNh5qMlcCx7QdjZPaJ6fPIKSWuB0qMbspB+S4Hebb3td
LIU/itjRlxh7z8NyuyURrvi6GAHZ4Sl26JlBrFHYPTeizCmuAJAKCQl5L+BbaL1X
xtJiw5Vin12fi+y1lS9NtGjsEfSfAYPBZOeaYXN5KtdtTpzwUC2+xN3Sxe5Heu2s
hhVPk4HwujDFBlljJZTEPaKRmU771aDnm8ofUeVMENi9G6x7Oj4eRdgq+etR2jh5
oHUY56BGdz0YBUC4K0kUQMiQeUre9FCTmSIpdOXLmOxR4w2+70wAXg5C03vY+cku
L9kYmoVZRIkQaK9254hMVp626RhZvgnyN57+oYWlU0/Zmz5c1UDUVMEraK0QN/GM
K4uebXT7Yabh7EcDwK1dLxyvV5kdin5b6D5rDHa6HyErmqE8rce0meYhA74XLcQS
pTCuDfmMr6yqntArxoQxAEggjQPALJ+tTqsmPfvBadx/7llUPrmnYdYcdwrnp1ed
B/l0/3vo66YpBMFm/QbILukwhxRWUTd03BO0xd9uSvlEreYSbtFiUYG3LdyiL7yr
by3V5XizOkA0AiGCpnKyfswav4X6RK67KufR7Wi6qZVb6cZ/ukho9wlpMaZ9OVfl
luxqj0fKzcfw21ymOS0PVT95Ck++cH45olapw0VjCnFPswXLnAONExlo3Welnfpe
C8yxI7FHsqVS+H67hZ4UBeuvXSwsu+9G/6vvdz7tQPCtXzoS+dYht7ZeC7YJsf0K
PUagSUs1kYn9lqSUHJNwpZdodCUDMnFpLnPgffaB/Oc/u390rDxhs8b1aALASNwn
xsUUX7kppyql6zfD7NEdCT0riy2PFpht13ZD2G0Lz8ceX9941vCmcHBU7Fk5wcer
l6Z9+S2UIXwowgcykdU9gnkSAb+eDBLc25HfpssEwIZ6j/wnj8J+MvSJxlrFt5Tu
XDx6/O0sfwOPBN8TwI/vBN+dVsEfIP4UZWpvkXiVVglB9yemc1zJryrmB9mhrwSN
8SQvILOV8zMvEmhBUsd/1SiwKPVXyoo+xDJ2BWLRL3t+ovuG+HoKOQrAISzns84N
hp3Sp+dLbXWy0rzSnKx/UMsTxbxfggH4aEGlvPFeUEpITK95IbwVaGRLZUx5FeZa
z/GS3/slgLw/OXd47bh/q7Daab2uI09IT075Uuyjtqbv7kuIHSVUyEcGvFHlVCVM
DUmiyUJDaeg2/z5lLp9UelnkiftrL1KfxbVrzx35J0xsVpCNayU4fIa9gVnWtjC9
B9MdUiJ8RXtAC4GETLHf5kv7oA+BvkIkgsLuPyThlnkReSYMGZlgBZTzeoDrm+S7
G0/ivKJeLrplmBHQxHzMJI86RGMffgeKOwnCUqiTHs4tA5TFBQPW5MPJ47IRzIyD
GcHGH7f5BvG+kb60Ruoq8iFWav8pyhmfyp5Vd+WXco4/19zTh9E2hlqGvc54M+09
IQdQxihBfq+m4KO2tzU1aNYzEYJzVs/LRQFRpUPvxRsdxcsXuApLlxgzfPSK3M+J
nf27e22Qyk2s6H0i78Lt4VSiuLEwaeDk8arjhxngE6fLwbq9z+oADk02qXR0ndd4
5w+G8hYRR7wwHCX20kLYqEPP+9mQjWxrUcGfwtv77BAPbs9MCuNPj565Rb6zhn42
wTyGQfGXOuAArklFqRtHLLYfQrfBtrNSRX17/FHBcpieidbg2TcvAGUAzLhMWZxS
MkyaZnZIhW1LYvhAIdmJJkV68/tp53Zg0ZjXRcBLTGwpEcEdSIxsRA+4/jxNZDry
oCNXSm8cQwZzLMgxS3WawGqRwug6q5qL56Z8jzcW7LlxOCFdLB1ilrj1vhLsIuzZ
PhYZ/QaUwkMlwu41NFCr+Wyh/hhJh5OMu7Vsa0StvT8w/UJ9AAVE764Fk9CYzujX
TZ1Hi8zwpMHf49Zg1QR9Q2YqMLhCmFssgnXfDtOn+cjKS1heyc7dij1TdbZJgQUc
YxzHu+JK+PQhZ/6E5hCigvTn/R7K2IoWucCBdp6MZHwD+e8mHrG0gpSjW4ZS7FrI
sCWATUIsnCNReKRIGztjx+p2BIWQivBfNzjFHncH6UdyVlhmg2o+gykbvTN6xRGR
cIRKz2cUYkVbCvdJmYRBIosysh6TnfFHV6wc8v2h7Q+WopZOwj3LBw05s5SuSuxe
DTv9lBhKUvcdngMAw5ybSg8p/NEhgNHorU/EsNPviXJRqpC4HYVcSf20a1e2E/7y
WpQEwhbUnK2bEQ7cK1dLgLG6SJeDqRvQ07n55GQiL1JsIImsJrTtVgZT5iLSscxn
tw25mHp46IGYOaLezh9hgWb8udA4hFxTekqOkzt/ea6wXpOMrQbLvOeIU5mM/WEl
fsZKKSqKNRrsRmRXwjufuFzlXS1KWBmpkDz2Ra8cCaQDsmcPhaJe6vVqhKZvwCQh
Lejb3v9GAJ20XfccSACQuHMaGUNG/b38zd0gBXNJnUQ7vuvaK5pjypgEkZ4atEzh
V/T1f18nxjMEF7wYnCfV+9dZF9PCAYQ7ZGfXwOwQMDPIxZCfEFv+5Hg3HQkiLWye
zVAz0rQWcCMgBUnf3rxSClq+Jk5JMesxqA7zUrMh+cUeFrz2DnhgDPX4emgIog9k
iCXbQcKH7eMCtvJYJd7sBWoRKG+oZw8kAIbCNokk5uxQUO74tcduqBdAJ1NS7H3r
W6EwmGYRZBlRF0L+ab95LHLbeteYRvdyCtCudHtKOykItJLvuJ2KYrnIW6Stv1bj
pWrSydTfpyF+bAk0o/osE4odGUPQYrzaCqYetIuqQZ3XXDtCJhJecH3KzZhIikFb
yZiTXgvAC6seJRE3zxVdHJPVlfWoXALOpnXyAJ43VrsvuQvIHpHlnHaCGzaFU05S
2CwfT/gOJ179Efw/vRtxv2qrIOPLwZClZ0N1vdEJPLLJWMXGen42ZSL/aib//6bW
zzDMwRpLlAIAQidk7oaFpZ5CvhpL0OVucV2iCYdIIBnjFJIGApi/Acg5FGXc3w1v
5n+t0/6o1T+h1rmmR4f56CrdfqXBLi5EOc43Fr312yG7HLQJnMwgJcNzvvCt/jXA
HYaeJjRkXblmKGfwG8jDp2P3YVgeYc/BC3t9gDY02pdwSS6AjTACo98wSCfDVXQf
qfEsE6HFvhDWoD5/oBpWQWdByGjZE6SWPOMdpVIlIBvgC7baKZ4YsXfjD3oAcn1U
bJoug/u4/EfDpwgECngLJKqokGMitg2PdsttxZyrPO/rybIxCPJhg5HrjgrLW3VN
dmALGR1XXAoAQpP1+Hc4ddtG+U92aW3U0BmPQLd+0NR7Oi7ZU/APcpHuV2/ELGpV
xaHKuyYa0qIM1U3X73UamY2jjh5798/ABLBW3Os3sZFCaTpgxU/4YTJ9Y1sjtKnD
DeBomk4WSEHyXL9HIx9k8TOhd9uTyPFKKLla6N6sx9XkmccovMqOGLMZCu6AhSd7
ybqkp6lOKwMKRCg3Gi54GRFViHLLGRX4fNvY9K59WbkonwOB4/RCc7iLWps8d0pe
ZnULSxZOMhKMO0T6lmKsb78RpNF4gTZ9pWfEco5JvfaM6MCNLguYitca+JThRnVa
kPLhJdbdvYPzD8i2Fzo/o/v4eAPocJb1aWXvYyONsRXBHAzOSKDvmdU6if41vmQF
rJnITQM7rl3MApzOClN1pG+E2mB+txj0y+GwMMHktUic+uAZOQd7b0m+na4FOSa7
WGctK/85WJNdHkYumE8NPDiF01JrTBLQyqLRsWA+6+v1dKdGrGgj+2ijB1yktP2R
Hj1IxYly+TRSd2QapG1zylAbDzygT/yjg4qSaI6eZz4mwQUDRIEn2HsaIHS8Y2N7
lQdr+5NPGyKPxrmc19KuD4T2kVDbN+hYIArDeQKBo2eBNupSWOnmKp5IWY7Mu7IL
s4P/viAkr/p0Js3R5rD7wOjgj7/shezG18p7aGkmRTM22ej4kvV8y5fV9lDfd32+
+hRdrD0sCKWn61ezR1yOyb0a+uXic2FSc+7oAOMLfHCo9a7Db37gAHEbcICv7R+X
odlsZFCVNQH+EYJS5p5P0Uam8kLxNeZ5NKj1OrK7MjPm6s1LGT2tknlZ7qEKZgrK
NrQWP7X9k6SIlzonAnJ739PM8A0hrE62HkSbNECCx8yShKPiisYitKNBQ512PYyw
CxtGM9EbsPKRMZK/0jLrihnTqComhqQERUx01nXAfPjB4oa9ItlFYGjHq/jtOZIL
nDBZiEpTltywR4XY7ZpuLg9uRhcIhTkJdyUhhOuuBWFKr5E9AdRVkluT4zwJd1R+
i6ueYfR2hFbl8Go09zF78xS7TNV2OHApuKnvN4Kx8UvoGrsZqzba/X9pPEs4kXMv
7Tcv/Cr1DCxrTrzrkPXVh8OaUO8HCb/txUybZgDf9ANSaaAsL9/STaL1GDE1Bvfb
D2AJc1RNeHf++AUQZB7uRBYT+Pohs9Iwa/Gw52Y6q0F8muSpmDPf0Lx7qQZ5SEUw
I6PWqMWHOP+elaunAAw6B1q8DGKjF6aS7AA8fl40Qup00EqS9Elt8uP/I+J6X2p3
rWn85cIMeQUb7w4NPxxtKn1bGLQWnQ1/Oj9qUV533m296FMRr9sGbnGe9+gwYvW3
UWLoJrsdyJj6AWyGHmTS4GseawOqtUDU+sxIyLlKCvgroxL/pFDI0iG1DLU67dlf
3pCX/nVo91MXzMuuTnsCBo0P8+G8y/ZNOR4jrqip95xlY5PInbiPjn45PPy38JIl
/0/nUFJ4c0dS5V75I6TDFirf2rmryZoPFp3qPLap33Ui+7j9teVFuvtSPMgPuEp2
Ft1LmBsUGE/9YbfWPaWAWYPnVKCDeinAf6NMdGOX9lc/uZJu8Q/l5wvY+wcjCRpL
LD3+tCxYWLQ3nNrrf6ODshKUewabFsVf9MlSlwOW1UImbdpLLTliHyE9zzL6QxoI
3QBXyN4tDi55YfmxChh4KWnoSuQHnswBazfdtN+fbm+su8uIv3m+/WO4fNa586ol
t74eYvoMgQ7gZoxewoi/L2/HXHLfRHTS0OjOkHabCuofXrRXJ+ou7zr5sqdJMSOp
35O6iPM7bHFmJrBWC736jDhC4d5S2Xu8VV3mgs7WcVgobPKQvPjRSzd4QwTOrUwp
jA9qqD3mZAoWlwZVhpRdEzWIttK08l+EdcLxSXDtRbhiRcKwkoeLcOMRsNgJwX+K
AzxWIO+4QlG02ij6Gs7Cuay+07ImH3jO02W3KGE4vkXWBKtzVI1MG/GmBmrRyJrm
UucEcuX4O5/UrrNLMdvFk5M2MvnRanU0urXgL1MR7Y0V3CaS3t7aXUO8s+TOuFuk
3Ey9i41b8mN3mIxjBxfsdacX9ZopWZ81uajGW8UumfmKh7p4kIYUtF98dt+4anTL
bdb+i8fK5sYeWYoVp7xIpZHARUsxRbZYjTehtQIzRHBidjsHdcNchIQfC4j1dfFd
gs3KuioEZSX1v+DIF29bUrirGoQgVGILjBNQKWjjuhSL0wA9O47TCNm36pRiZxTY
00CpxOsiyk0mU+Au1RYSva2i4/EO1jFfm1k1YxMPZLQXfa5wpYnXp20pbsRJ4ZE8
bIebxxucRYCX4DXhw/f2Yx+UiHZEveEwmmHVTigzUCysjORL5+qjIBTJUiHUDzNv
gGtBsuSVHJ13oaF797m6QMII88OXn0kayYNf75pzqR32ZVjM47heyn/Z2n/NjHu6
fZJf8nDRbecIJVx1fznoy81g9b6L+4bj2tK0dN9kcAG5en+1jaDertU9NiKZapCc
cwH/EaTBpMtSMGofA9JfHsLoE4lPLbujGAoGOXAsOefNGVQgxFfrafZjfi8DUPyW
DGTiYC1bvd15am6EqXU9xlGtOL+0drdGfh/0LvqIcKIeKqe+bimi0RguK5N5v7eR
Plq4vqhCiQxmAefBhdFdl1ioya1vcUc4nduqE0TDK1FPBuMBN4/oUX2bKSf8emnS
hxD9NKp8u0p1MJtjChrz2hrkvwKfD2kIgERNt2rB3ZNUIGKcm1tIB9xhSb3irI0Y
PskNguRMI/4t7U+ObVS4RbXkDSl2CBSBH28SjRfz2ceAl7C1OESpOS6zphbwbxSI
sh/3NkiiyjG7NPJHqcoXl7Xvig9r86rQdaMiUW2JY7mYn6u4N31zQVc+PVVBp8ak
ztOMUMPtecfUJQSzWp+8TQ1W9u8coFTCCjyxpi0TBXxCm5PRdERTn7WSDGj/qkwk
pJQLqt0kN0MtNabpchbbQf9cYXRve/HuQXby4agYY+Ka8gJeycdjVHwHOTX9m9fA
hGZGpFphmoitzoIHYpLqF+WsgO1Ty55S6n4X+B7fB5byaQuimVjapqaX9bGbR0Ko
c0CiXYsYL8o4oEz4kiejKDuBv+O4Q8hnmHx+sskML/lmMcNQPNZeJotbhFCXaedw
kcgijYGzYvqQGmP3Pj53HlDYS6rKl32p+rVuxsIqKuEx7mODr2wGe7z9PioJKKN/
fGa5k0Dl3bkUt8FwE8xXShcsYa8mcyAXY21U4keGSQqnnkZLfNtcd7keXwHTJAji
lZFo0Ar8pbgn/u5TPgg0rDZqQoHOQ5dCw+z//bzU5SDZ+JAgTNW6YEllPBP1Bkvv
5IVPdvm3Oe0ILQTfCVD41gaWvisiP6I/UDe0VEoLlyPgduzWCNpi3m6+tycahs97
bDXjzvb5kN2tbl7yKKIYQFFHyPwJqYlWl1yKX7Bk6H4MTmyV6Iq7zyiQUr07EZX2
2eSA1h3tC9WCfI+V7C7ZPwGwNdMPd5T5J00aUoNB0OirlO6athI32A9+FFo8zqjU
mGSOVxGZO53ExaR+sIxEILdT0W/TTfRvn0+NmHNMeub8heoDmpZiL3Oe/atEO58N
fU9ckqC/JFfSW1taxG0NyxP/nq/4y8ZBOiDgcbgFO+cdDSTEUusCVR5T0vYFZl3k
5SYeUfpAmG7XEHdjP3bRKVh1SzqelAmM9CFfEyOCgCYAAku5cGTZNAotyinm5wK3
h++6ur8wBeZ+OxIYe4sopt/0EhwBeEs5ztdJPaCNxwZJpo1qb7C9Sjjr+HqTSpnY
05y3+JyEkWOkVSW/haJSYOhdSdYLb3EiBFjxS475cnWFLSR+y0T/w6jPIdSfu8BL
me6xcGUC6Vdr7Uao2MWp938+J7HZcoNL4OeQIBBsU9//WNc4zG37TY77GUaH6kud
g9Q7841NQ9pNfPTrwxYSI+25AXGqNLd7cyVL/ZTMzYGd+27McDfvG1iIYtGEcvse
kjwOoJ8H0IMFRh3RKLpOIMKEusyMi/QiSXgIsaTKy9D2XkcbebDVUcOCSOGBPAFP
8kRhTHc+7vTTKENqE4HjhWqMKgL1fQ1419O3rtB/f0c6OWfKM6mxBb8SqNsP77TQ
VqmxiCYxQ5HkzlWypu+k3CA5c0nd4X5TwzG6IRgYT1/wMSxL01hLQvN/h7xmvbxw
Jz2g/8YFXnspMM5AXWhyqaCIZi9xwNeYo7RnoacYnrNVLRXOO3OlNDCQEAqq08IE
og6bSHWGeu7fLPrfv8LhDN6mkjmBvlQVWsY5acHyb2HE/DhGVjPplFarvh+Crp08
rpr9Em18h/BBVkhkTrDj5V+1or7DeAYa0pmOn6/A/68i0sh9ap9KNwDhFIFpr1Sy
o+2nAjtUYhryKL9BgcFuB2n/v5R4NshAUQ0Ht7BVx+CgqRvPDPeUA5cmP/yyQyOH
XmZQRfulI3DV5xJbTd/Qe6faF8+ymyJs5/uoF9+lL/A666jvGsTQZxtDVDwMqMQJ
y0MTis8NyShz/Rt57+o1V1DbBEKakembSx1F6Noz47Ae5+nibSjoACGJaLzlKyT/
ZZGETdpAucipw8xX+kGnPXhRoeC8IFuuEfhINv1sR/Bo99+Iwluor9prWP9xwNSK
gwdndqvp0Z6KyAkAHif+RkJdrfHT3mysOFJEHElQe5/P+rsrHPCyhaKlV6auTVQd
N/M5DWku0D3EH+umZeYFE7EML3/MU6YmkRMTgFRXaOxaPHyFA6xQttRnWB1GPE8D
8FMCJ1q524TF2OT9+6svCQT/jhyfgHsWKpb8AlgYuYXciVocqG7aostKUma6iGD3
Q0czCXXppqqa4oy5/IZkpah8GxUFxPxr5BZlfeqLYv3LHsWUjWKFKQNCNA86tOhH
BOhQr3oL/Atmcdm/vRuCOoXVllkPLRTdMiyf0xm4mQsoq/lzWW23S66hURTxkrub
/n/yrGmPYWpV34gOk5Pomtum96DJmLAd50W/0n6mhcNjTt+7xE7O8yAZXMMsb5Af
/Eumj7bem7p56JJgMlUA3y8U1cKFD7LjmTxE43bmVjJtZiN/aonKwwu1F+YQ4pFh
EU+7SP72CE7IwWKdI/L4HaA6qOA7AT5gldYjVhjSDPBNDxrxXFTzkaCVJuj8tK4e
bc2lwenBhdJEG1JJ5XsFGCyT/eMjBTcDhfqB2xv3Fc2Xt++stM1hKeJKgrRBCiVV
dNnVxiJPhXLx/CUdihOzbc3KIn+GVyBWpEiY9DOZvT75eOs6Yc7UY5mGaWyxnGnb
QrEtW7DyTMc0nKFYHXfqidbn+UVSEdS9/ABBnMrCP6uve1jgvgY580EGt8mc0b6A
BKUQTohHn9mmD4hvfbyav1cyWeFjWHg823/8n7qevTN9reaZkaAPHjAQOWDnMKN+
6cBS/dZAzyLaAJcf3yJExwUBBXpK8vIU+jLaUbOYkmUqyr6lXkTaGJ+C3sJmRpSC
tBFU1PqWNqyB8TR+FZlpr8HOcpE0OTP1plQCrIcCqJZfgXCIlRrq/v6Jnhr3x9Wz
s8fBSQrhMbvyzumbf/8FPb1MY4hnJ+qZY3VtZYnXh3X59QYNFt+xYNyMXD1HWZYM
D3i203UDbyTDnUUErAJkY3heK3E9Aw4Rl2bri/YNG4OkAwB8Zkg6z5L8gRQ7Ozol
5GbhqVtWCHtNQe2Y2tcOSt/tt/ueHTBOHeWc8HdauR08w42a3uW3YplTe3LTdDPq
WNqS7Z43UYVJt24wXo2VH11019+XGGMzmORbYxM7apQ3S1DspBwfsc43G3Fkg5Gn
My9egwTYWeuOUEwCRlz5qvETm2FK7Af/X/F8ej3kHY427J52lPu4SgH2+2J0g4cG
ZtpOSolAlxf65hNYtXw9LSlLM2G6qTbxJBGEOcBRf6rpt2YMUktu5ykgF92llOXf
bihqYPpgHValNi7Par1Sx7iHfdgv8B8UZHDIbB3pzTQfk3GQ+aZu2ZjQP61n+KC1
AY77FmRgL2PbU+UniF25xBB/VlklQx2q8AudfcuoPHAD2uBs/t4qBU+XMkdZVet1
OHatdhpZ3eaTLa46NI0icNzPO2KE39at/N8YpICf6PCIYJRuRDJKusNsmaNJb5YR
FJIsIQoW2S7UfJh9ED+m1EB32d2rEL0TrlxA224aoTp7435nQxUA6xjpFyicOUGi
GY4ld5CCtuSMFnxQXcftm9rjZ0BE9lUEpZh6tbZKTubtM9FdO+wub58PZPSaYOtd
ve0srJ0h8ghz27uh2+S9xttvm4tlbLnbSH3tIfTDyyZ326u/rc4zHCHFzY8e8pr7
yEucFziz4jYnsZhsPbT+9x+1a5RXfz8rhGGO5/Qu3tdc/WxzBgt8mv8X1DOroVWe
vqU4SCuZrvv6pUDUXWPYgUowIv4bvgU8kot6nxwaeyHUtdYJvd6++dhk28zXtMeW
Ner7vRauuRm+0x2JET9WmShG2TJUUQcD+vgitCKm20aoT131brRKx4Ug9Hx8a97c
JsYZz7a3JwQBtBpmegPVhkPKR9Op2FTFX4ARbnNDTdOxFd0EovmTNdN8Iru6cccN
hQ6i5CaLJxvi20zVB1ObjTLHCs7m1sC1noxxT9cokwEm7F07iEXqedbug1ZXaDnJ
fsXfd8xCVkdtYw5bckIcCj5ttsMcirIyMNGu1LJRwkmtpaimVQ03s4EiRy4C5eYr
uGKZTAeJzgrDPQQtUT6cU2i1pF84F0Og00f9EFEsGQUu+rQTBdApBxutQq7Rd9LY
iz9syyzaiisUjwpU2tmaNBPV2llRhSZjEFdviEXRne5F9mdGRszWVpQLVmq4k2fM
0LQWa2he0D8goIzXyBKlkMJ4PwTyjjyoiFgi2/bbk5g2jJlGNP83MYZ89bY+I+DY
ELpOeDm3VS04zLsZn5Dr4V8Si9y6gfgc8ukiZcwuPUdacxjQOtfJG8AZt+k4ohyV
9RULVs8wwuwHcBuZByr6YU0SKaXuP/ebOIkoVXo4eDFHdopPkJaUEKvXiUCos0Q3
7jGzSjtZPV+EkFE8rkHf7LBqJrJYPVRukSRrYPrvUmBCQSQ4AsbuIQUbBq6Hmz9B
CX+h20kDzh08qGmRkgSU49Z2Sri6OnkRla2Il6YVIer2GHcSpz8iowUnakv8KVbf
nJMNEdYWdJVi8MWAx5I/4i4YrHK3GhR1u4re7i4lERcmO7ZVsvXsM/t9xriq/6ew
x5ajWlJxcwK31PqQtcd/+aU68x1DVPKHxx6vKXwxajZfDRfK+keV3FJmKuuFa2MF
k+GmJb+21dLtDOdamaAk+K8lKoZJPOqBCc9ig32pHnYgBCY6wTwVqyNJIEP9yGda
4pGERC/HIvxUjhjX+ft3aR4WIK3iCrkyqZDhAECZ2OvZdgd6l/VuIdCxScRc8flz
Gp9uc2MeMWERTAkErrATvQBoY4Rd4ktISXsnicLULlDWApfOpuRJa8CJMfr1Jjhh
2J6IDtb/GVOjJs4vDHEEj7A/dXV3R9B4MjVNpVyQ6ukLUPzglzgEtuI97jEw2Bpr
as5Q3YuUTsOCIwJpgzShP9Dhtx6WAwxmdgowgiViBBBfpRXnRtydMWLVqrsJFS7A
MvL7Z/B6esHx9HfJQiXjJK38r4PwWiF2QlDmQu+bpmAnNB0gSAUGymyc4O1ku2MD
i0fSZ2zImPTWBHs1wTynt8y16hgt8xuBNnmfDJVxLRpEGgCHyJcm/zFFasKnRBQU
`pragma protect end_protected
