��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z���+4eTc�D��)\����Ķ��?I� �X��L�����	zBw�]7�^�������+�1��E��3�C?I�.�9�-F���PB��Z8�̂�L��>��W��t�ۯmS�k>F%����`��7�^�@c��P���a���>�[���O|ާ��/AkY�1ӫ�L҅��T���}7�	B.À�3� <Ns��>m4�<t��E5&��vU�BW��+NW��vU��r�஽�]��ݨN����R���kAܭ�\���y�� �����L0�xP�4��X�g�cm�N��s1Ʋ�2�&�VR"����;ظ�P☫B�v�o�;�9 ��~P��aw�����w�6|���~��`F4SP�	#a׎Ǥ��{��(�o��*(d��\�n�� �b ���T�V��\�`�w+ӆ'�b8������:��#��	w�t 7�H݈`ƌB@ �%4�I=��bKE��}�v>M��3̾�,��-���:�P�7��qeӉ
�N�4�-X]<�8�-��_�ޅ4'Ѱ3^�l�_�a���>�\ʵ���&�v#��d�{�i���+�]r(���[�4����,��Gpz��w��Y�&;�cˎB���P>ri���c|����f΋e����_G"x{�R���C�=&q2�tE
,c�h��ɸ�At����|����t�����LPN�Կy-��oI
��M���A�sT�񼏨�]�k���=��FmO�(����_�!(e},�SG/�Q����7�ZI�����C2����CqN|V1�v�\�4OI������3�����xO�PdgKg[��Ր���3�+�!���V��s�&(��@r<hՋf�V�(X���\ț��/}��F�Ek��	kyC��G1�S猭JQ.I�ۙ^�7\�G�o�Uc��/�M�O���}\8?�E���§�����\�`��/)�څ�W��tt����Dk��
����?-��S�>B:�Zo�|Q�v����C�^�<�@�Q�S���B�󐕧ҕ�MPO'��P�T���: 7\�Of���7u�5��(�����(����}p�Y����V�����2~�G��8�n�[�ǒ����hJĖG:I*�/�u�@�+Akk��F�c�+�/�"��@ZP�v}���?��" m������l�w_Q͇;چ9�k�x�*I��4�[��D<�;l�kva��1�d5_�bm ��U���ވU:45Ks��/��J �Kz1���C4�[+�I��g.Zx�"˶sez��bӴҿͮY�����'�9X����7h��y��6"��Kn�O���mòþ$���i���ɡ��}�v�vc�˺$���91�/���^ܫ�{!'���r,b�J���椒u��^��I�\R��{�\�~?'Q�a�pBӒ��O�2"E�G����������G�}-��`�7Ԧh���σd����r�N�N��zi3c��׈e����X& ��4"(�#�b%�o���,��[�`�J�ׄ�����Yr�6Ѩ$�y0�����O$? �(�"��[e���;�֩�w�����G;��`R��{�i]���l�y��^�ga���ss�6��&��+�Xuw�mdb$5�0 ͩ 2���=�0e�&�!���f��<�o{A̋�c��ʺ���ݏvx�0t��Z{����l����(����.K����<����6�{�I3.d��jbv��+b0�pF����?�鱓� �o�7��4��*�zњ;�ҵ��_7�Ky�٘<�l�F��~�¿/�hb�Sb��&��������W=��Ӽ��ϙ���6�=�(%���%�<����HW�M� �P�L��.HCI���j�UȒ�^a�K�� ��&|�q�o"C��u�/T ��Dv���ϲ�&%@��<6��k,���N�p������L{1��* ;&+���3�4� ׺��,
�-J��sT�����\P��5�(���|O0�9J\��5$��Ȃ�R�CʌF�0u�xPN4����y���`�����/���N��g��g�6� ��-������k]u��`T���ޚ�?��}��Bd�-5�C#@�`���Uv�V�h	;'+:��8�vm��O���M��7�FMd���ib�z�#��/,åf����D�� ۠�=d.�F�T�Z$�j����0�,�-�`��!�ɠ�T�N��q�;`L^OA�?�*����$��.ζvEbM���^���"a~4�n��"��ۚ	U���tI}g�c�2�+��Cg�s�7s���Ĭڊ+ir�����Sdv�v�`yF��y3c�Dc_f���N�H��6Ur�ҫ�l�U�Ȫ0����8i��p���4~.A^,�Km�[��mr��^��֐��,@rbMi�V7 ��D4�C��W"c;�j`AJZ_8�h'���{������e峼p��l�4��x���&�:���uV�~�<޽�����M#H8��I��U.�r:Xs]�m�������T:�fS���C9�``�3�5�^<��c���?�\�}��0��~�Z�L06�����~r���ȟ�6c�[�²O����bV�� _A�tu��s���o �)ġ~���S0|sr��m��EB 1��p@)	��͹��3�	�;�(��6C����G��"�Ί5�f�J}7��޲+t��ydQş/�e���~|{쪧
3yϽ���Ƹ���[ʂ=��[�E»��T�~'�I
��3��DKߦ�O,�R����F����`-9��tS�D�C-���sUM8Ƕ!i<�5>KW�t��7Y�Hw���2__V�qA��,���c�k�@s �_#�nF�ثiԄǧ��⳸�9V
ϖw0�VF.o��u����͵_T�g}���2������)��:��TB���G�g@)Tvs4T��W��cc�ȧ{�(�=�5G	B���������͇M�0��#t��\r��L������y��/Aڄp�(ˈ@�QN9�1(���ʕi}�L����i�DE���? �h���D�2,1CRG!�(�ɜ(�7H��}�u�z��s����&eA�H���Ӻb�i��֦|�+3����$��W%s��ß� ��[�ζ z��!���[ܟ��@�7iy��~��6�l�\�O�j�P�6^��8Ē�f$2/�
�,�Iq��E��h�:+5�9�������=���\�1���0��0���ٍ�.z�,T��c9��2�'��ԑ����c�a�@L�u�^���0�S*�[}�E�3e����t�:0Q�N�ĥO ��m���G�����]�>�5�����-�7���@����~�]Be�����6W��	Lt,%�?V�a�e����<��-�l�V��~��NPn����[��W_�)Z�=��v�������T�5���ǎ�=��`�;I���K7��Ҙ��愑FIG����OըN�����l�k����<� V��=�S1�Z�cT.����1i���z���,��\�\�?�$��=�w� ��W!X�L�J��|��3��j/KNUFl�UZ����[�$����BNV��{�θM���n�	�B�^�˷�|}k��q�)��`1���6V��d���uX��W��" X%��ej�f������!,+Q!Ke�'W�N�T~�`<�B�Q�+v �Bǝ��++E
����W ^Z�=Ĭ��O"��P�/3�7�M?g$��Z�3G	W���@�^�G��L����}n��|6n��~��5k`�y�-�2Y�<K��RA���I�odk|	�l��C�R6���]�b��, o*O�opt@y��se&.,g~�����x����eZe,�W��ʺ�H�p&�霛FT��~<(��ՑB���X�"<���U�f��"���=f��=&b�DUܬ@hXJZ�_������J��|m_�М�w�5��ޤn~x��g,N�����㲅�����E��R��+G\3�D@����="�@�ĥ�J�rm(�*j1#a���h]g�خjƙ��T>σ�;��%�bt8�|v�[m
�E�G�l;Oו�,�(�}�^O"�)H���W���SfM�t����"�heih:�D6�;J 
�yx�9f	Y<�.����r�+bxg������*������s������L���'r��� ٺ��Uʎ?a�t9e&��"QRm�7ݨ��v�n�LZ`-�ʶ-ᐕ�L��[��I��R��_	*I}`*�v��Zb��~��-mH97�,͎ja�R�7��6w�LzW��?�Ħ�5H��0]b�y�Rn]��������ʡi�6:T%�b�N+���s�g�%�X�TuL��?v��w�WfsED���� ٢������[�~��8j���i������#�̉�h,�L�DS>_^�ը�ݳ�$����������M�znD$��{˵*�,� �BkJ�`)�6I����M^��>5`T>h*+���8�=�a�Oy�j�5�H�+���*�0>'ʉR1�Sw��V�lqo�&�(ʀvTU�E@�O�S.���D���ړken��]|"$�hK�z������ƩnO7[d�d�΃#e9���^
�{��'�sQ�$�-��.�̤	8Z�8�dʃ[ۂ�>vam~:��?�.zCd�m�Bq���3b��J��[����;�|1`�s �*
9�pГ�o�	��,�D6�͗M�vE�f�(h�%��zMH��^AV$�{&�i�	b6)G�
ݓ�3(�C²Q���B�J&i=S��;��̏T������N�BmN{�tV�A�JR��j0�B�&�ُݻ[�}����n�@kq�R���S�ٺ�)�m�%�*bvTI�����(�蝧�D¿U\'m�n&ߐzS6-��(W!\��	����|1�v^��!V�2,���u/C�� ��R�;��k��`�.�2N,��|�w��>E���O�H�pC�'~#�?e6�,l���(�hOHY�tx�~-���^ء^�󧉵��ٺ��I�Ge�w��v��)��L���%Lt��4����R$�c�0$�����%�%k�ڈ������o�TZVX&�~=p�;pL��v�ubI��K\�k�XY��G��1�)l��&qw���ً��J8(N�����.d�]�wS��"CpqLd��� �:��pg��y��މaěl%݂v������t�(N��l���1R������6tu���)U��k�Q�	ǿUe�j��y`c�\�L�%N��*CQ��[o��G���A3�J2P�2'a=1# �Q�Ԥ���1Nl:ҷ�VO�Yvr�̅{�)�S���;a������y����414�Q]
w�'&�z+(b��Q��!�3s�%IQZ_���L����J���%v��Ζ��®k�<'����w8�D��w�󑓬�DR����<#0���b_���!Q�l����s'��Q��΁�[4IJ��pk�z�m�tGq����id��s�I�Ҏ5@���`�/���d�(A,�&ɜM����e��0μ���łT:S�N�:���~�v�343����$x�a�P���W@��k�nI"O��bdF���Z���6ٌ�[U��ob����Q���7�j*0� �㱱W.:3'L��~��;�*�,�v��~	cE�8X�N�	���2��kF�9�yV��n ���(*j��j��o�5���~�	�d�F��T(��jkݵj����!�!攱��4FA�������g�m3l�W�+��ہ#r��$Z�/���[TJ�k���X���LT�5�	擙��
�Ggv��kK�F
��Liٷq��q�bCB�	�r^����N�-��άKUy�K����L