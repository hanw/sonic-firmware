��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z�)�ŋ��6������}?��mK�x�-��痳�6��3g�w&5�pb��	�y�1�� �~Ї�ԏQ����*dMX����H��	�S֋}W�K Q�"�z�4r:�X"��=���L1f��,�$��[8� �M ަEi^��u�33_	�C<*���:��b"z9+��M�*
�̀^�
�銫�U�\�м���O��#]܅��
�^�}2�1��<��2,���a����t:�%b�*Z��3��t�ٽ�;���2�]HT��(�,���e�HAA�O]O��E��!���&0�S���,��W�.�j��${��*	�R�i�V�
������xȎl���ET��`G�����¾j@W����YR9��bf�T���(�[I)鲋��,���$���϶q�S�w	�b��xTNH�vc�M_d�Ơ�z����يd�(�&�v_bj�\�,���1���S�\d��y�2j����\�' K�]a�A�
�Gm{��#,������C���<Ŭ�5�;�3+�1�B�i�(�6��!,�qj`1�n��#ä
��d�ޕ��9�}���Kc�c���B���'8�:�aY��$v���UdX��fU��`�8;.l~Z��׽�H�_���j����?/e{�������f2v��c��j �`(��Eu���Z�Ļ�^`�	 0Q�?�/:Q�������cv u`L�;n�Z�t��t�Ț}� mN�p-K���k�~g��i;@�������C rE69u�+�$aZ�N�+�s:#�o��:DˑJ��x}�#ɚ�`[Hc�q5�[�M�b��� m��=�̣D�����Rg�Z��[�H�ヺ��s��e��:E�,�A�}����+�0�!!,��S$f�Ydt/�0c���MFx�s���L���X�_�b�RGY�"m$j�תh�}	�����Y���:��������%�0��$�E3[=]0�L}���IC�>���U���P�����B
�������(y��K{����+�,�h>VT����Cy�(�~���>����0!�����$��*���&�a��^v���N-2�h��&������R)'
���7:q���b�W(�7KV 0��mdH&o��EKu��l�2q�,�л���翝�U�_Nb�m�x��j�*��u���=�M�L -@�Y̺Nl�NS�w��_\ �!G�}���ZX@���V�9��A�_�[�O��jԉ���j�+.u�/�SK�mW,'PDc���%j�|�M㏢�kl10D���,/�x`�w/R��ڏ(�y�� ]�=e�e2�p�`^�п�Dk�u<��9�%�,rP�m�k��{ڇ�#���_O��#D�����O��a��Ґl�l�=R6��P�z��հ�m�FJN��'�.�2Cc��=�� *��tV'�7)@�@��u݉�Z�$g�Iu�e8e��&dg�.2�K�5�t�2C� �f�������;q�he��"hS`�Iwۮ��C�=υ�?CR��N@ޛ���ԭ����5��k;�I���㣰Э�5�%Dv������8�p�2|���z�FY��ʕ��̞��h�T�U�E� ��?��l�B L��`��`�υ��Q�$������E����>�S�+���z���\��W��=Hr��˔^f+S��J��p���<*a���gML��4�`�c	�n���~���h��7A���p�L����Oe��E΂����~]d�"{B�	�!V�`�=��a%���Q�1�s�%x���MLC���#�#�J=�ZRI�^V�j��� KS8{u��U�Q��^3�֐�
�
`�n�����iS��)��y���c�:A����U0���D@�%)m�|���o-�����ߧ%�c��}�$cQ��Јw��s��MP�ý%�C����6��*�}�â�taL���9�����K�$�h�䴉�LuG���ӵ��Z1&(0�I��A	��hC"%����!iwav�p���;k�Md��G��E�,y��r�T�B�W3a`I��?ٙj%��⩯�1���o5���m�?�)�$X�A�c�����&��T�K	��&g��O\+	ۍ��t�#�Iiqj�p���?!y��-��m��_=�{�������ܸ�)��#q����L�-�L���w ~4�x���O8���i%��Q�ں�6�l�+\� ���tGS���Gw\�=ZW�J*�L����9"��ߞ���@�ŧ#n�������`���_� 'ʄ�.�=����|	䓙ϳ��I{Gp�1��Y�7��ۯ(�uk��SM�j��Ј-���@9�Z���p�eb�a�ۊ�Ҹ��)���
&`�$�q3��T�[�i��(2�I��[�= ��,�y��(ι�d����y>c>���#]��$��Nsɝ���+���n�k�.p�KZU�t>EbI�¡���ڮL[�sY/&i�~���:�75n⸑��Z���ߋ� �aw:�=8��2�Bͯt��Iς�~X�:y�&�.*����?}a�*6��rh{�k��Zb9�
��&�,p��7^�ӭ���e�\ ������?�� �>ӡ{�z9��1�0��C8CY�����SU��:�k1w����w�d��F�޼�3����!&���gS #������U���[7� ��ܾ���Ѷ�m/��{���Wp}�R좒���7wߴ��Q�,��`���F���s�/����wBx�s�
�;������c��@��U�������F"&u^d*�����Oa@����w�p�ӝc{��S$�%��#��082��ݩ;�f�Y_�(�A�M��x<���j�,��g����c��i��_���}*tJ���Wg���AW2SN#�3�E������S��u���x��D�����c�f{`\�ڼ�1~�R9 ����� 4
��Җ�g؍�d����E�+<O@N��Q%��9��7��3hCR�J��73H����8/�ǌmy�����Q���5n���{�5�p�e�J��)�S"E[�' ��*�B�x����[���0@2��,l^��k��Z�2��Q��Ⱦ�4�������b��|x8x�7'S F�������jf('3}F��+b��U���j��j�bÌgj��E�$ذ�������JU,��+��ԫ��L�Iͬ��
�"�D��՗Z�ô~b����Q$U������vR���葝V��	_/�#��� ̸p��/::<D��G���᷒���?55P|�d����=��������Dj��c�4�ˇ�d�g������y3zI��$��mɣ��U���-AJ�����X7-X9�LmQ�0�9i��V���_��%����<��7
4��͇�7s�>�vJ_����$��x�-���&��8�L��;��񲀃e����c���8�6~��tzkϾ���y�%�ޏ�T��