��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z�V����u:0��,Lk��?.��p���� #0�]J(�_�"�$�K]�wK�Á�yU��_wG��{���0���jOGM~3Σ�����l�_�Ɣ����P�sQ�&av<��TQ��=�;�.��j�M���4�#� :��n�G!-����p*�6�7����˖"Oa�U���˦���:U���s|����;�O��������EQer�#X3l=��_����|!h��߀��>%9,�7]��$E���hcu�&����u�1�"�M�G�pW������w������O
*��)C��5��t4���H!���m�΀�/��lO��A�+K�:�+�V��8m��j�ҙ������K���D�i�޸�{]E��Y��{�B ktm��6��D�"{��&�օY074r��ICv��"�d�iڢ�6��0�����v����9�^�^w|�ϋm�G8.Ir�\o6�iD)�cm��׈����iK���8D��|C�����H�fw_�6��zz6�
Du/��؏bC�+ƍE���t�OyT
�iI1��ȋ��m�c������T�N�e��o����}X
�X�;VJ���"�����$b-Pg���D�M����%b��J�NC�&fC����+?��}�Q�j+�a���K69 
6-��zIlO�5������)G �,۵�ofJ3�H�P;�����/ӡSO�M���1d���ʆ�����lр�t�*�'�)ҞK����r(焀݈4��G1���M��@J��O�2�2�0V'�,�>�KuT�+��a�|s5K֠uk�a]�]1fd|�k�پ<�<�I"��e�A=���/D�m�����z����M�6��8�G��a�?%��r�E��%�u�r���CS�*��J��Bx7prjn���,ZW�K�a���-���B�������Gp��mMܫ�>�w�fE��Cb@EuҶ������C@}�|����e����SV�����[	����f���D�.����{m�G��@AN��P�uԶV~s����$������I�exm+���������/���pڀc	/�l{�\�1j!t�X���qw`qX����le&?�r7uٚɯcAm�����ԗig[��_Q8ݙk��9HcB�a?U�5�<ϑ�1�3�����5GE8�,h-�N)C7��
����u4j��j%�g�*SN43u �z�J�JO��z�FҼ$B���h8˲�Bn�H&?į	J<��'�:��.;�R��J�N�R4. �·N��2���Z�>��a$'L����>$R!��Mc���:!��au{�(V�x:�1�?���v�^ݣq��b̓bV��Cd����Tz[�D�*���qev���55�������%�_��ɲ��-2��ܸ�3�Wln�{�!�e��j���5@���T���Eji���x�-6y��h��75i���P|�W`�NI�q}�ΫӠ|R���ʢ�fƙ ��Bɏ���\��VO!_� �ާQ"'�Hq�-3��_��k�p
*�3A�lfD�lX�*"����������DRX��e�!J46kKVM���k0'>��lTu����
���'��H˱<�z.}d������V�\ľ�Ƭ���d<�����}^��%��;��������`�݀��>a��'��/��ʺr�᡾\��z����Ϊ�J: ���M�n�L�?a��;ִ��G㶱g���u�B�]<�/��%��d��9�m�r���X�K��qjnfC�h#&fM].e+�:�����Qr����cٕ*��zG<{sS��N����X� �F�편����E���}��q9�S;(��;����rm����+�����#�4��5�(�'�ܧ�J�./����ci���[�w���W+[��@S�$]�2�y����#�9����Yÿ��T�1��TlӨ�٧�1����l]sh� k�t):[�������1ݙ���n*w�F�ev3�b�,�ҽ�q2�}�	+Q��z������PXh{bVkrw�j���#2��8�|���Oh�;��zڸdŋ���ƒ]&0�h�������7`�z�K&zc��d��S>:�C��O-���e'��n�K���s�%����y�Ѧ��Qgz����csگ؋��(��p�1��,�`�I���L
O��QL2u9�|J��4�x����d�3�B_"����>�1�C�#��3�ػ�##) q�4xN��Pz��x��i�W�����~)��4����b��x�0�������5E7�<^��-��.�<Q"��uP��z�0�-G(O�AZ�qi3>���%rd{5�""jړ2Ħ�*�3�q� ��E��T�e��B��=�{�G�.�<؟В;�+}�^^��wqrĠ�w��yU�Q���B��#;띏|j�B�Tiʶu
���
�߮(�.��<��`aꩋ&e���>�3��lb�*�e����=度��tz�ɺɽb���b�_w�}��!z4g1r����-hf���9�r��m��G٫8N�v�O����0B��#k�W�1M�>Y�,9�~�b��[�u(tz�
!㗯m���-�"���D�I�W�$`a�9���Y���h	SrqQ�A����^�ÿ�O��3)����h2��p�>T>Tl��*�����DA��B�X��M"��}5>+�@��<�Р�9����ΤR��3&(��=͙4�\�J&`�(_�k���	m�oz�')����OZ
=CCǩ9����WSm���]Jt�S^��`u)�����G%���ɽԦY�'
��rS��uL@jv]���b\�٢PAZ�P��J�5���A���2&��yN1:4��ۻU����4��k<\?�%��s�`c��/�e��biK�=6��A�6��7?�a�E)��[F�s�,��4?�5�eFl�x�Ubb2�x0�؈d�F��w}��ǿ\B�f�S�ވ5�M�aM>�,z%g���5�U�:��!t�-��EQ�|�:{e���X&\[��Vl+Qڋ"oI����dϱ;�������#G1�<+��:�L����ϿMr��b���Ș�k�z�E��6�VУ�⨮׫��<8�`-p/�t�rR����Gvg"w��&�����Q�S�O�֒�F�i���앸?��x�V1F=��o�f�=�˘�D.)�oǐ_��]/�
�(g��{��O�k4w�w#eA�r76��plA�ؼݱ����h9ގ�7ѥ[xA�{���L�D�����SW� ��'>�0֣�8N$����C���|�e=>(�/��VI�J��
���D��Q��T�&�\\	�	bfy��ޛi�Q��h�,�RC��"�5}��<Jŉ��>�X���	T��l-��b�%OX�fU[
��竵��Ձ4b�%7�v��J�.�Yί�T6tmW� ���~���67��~g��x���G�`��@E��s���%���ŵ�T�������`�?���RR� Չu��V̹��NH�f�a�yܮV� Q��T:� m�/����aR3�0l��Xg �l�J����w���ǋ���˂� Tܑ�b�yP���J7Ԗ�wK���$��4�nQӪo}R���|��t|Ef��@VڍpOjj�(�{j/RU�a��K���6J�8�P	��"��C�s(.:k��!�J%�l�p���yo����z|ԍK�JC{ݶ�7&|�̓sZ�6��E"S�?