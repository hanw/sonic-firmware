// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nWVwbdqsGtfpRrlVSxeqM7Q3zAmJ5USdmwGSBS8wXozVMgKSSEWwk/DqflbhAyRR
5RRdm6dG13D+U/EqkK/FRjkXEiPzZ6JmqoiIwaUJTqvL2tMFqSficrT9SmeTb+zI
z5w7tZ/NDIzRpVQ9Hj8MvLLKZpVLd4ZjkIconcMAZSI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18864)
uJCT7y4K76QPjbwhvFw1HW3VsTtnH3e3fLcH8WwsveifGXJiMR/kvoPIITxAF3g+
iHgefF7jvOKyp7rVidOYEj73nR4GwKesNqD2TprUbLqQMC2SBx2Pm6npRBZJSKmU
LB7alIc2vZ90i19zZ0kj9yN7Sg4/GPErOc6ywJt4Hqid0yOTKWV+llOMOhO6FN+4
qeuVEcPrFGsWa03V4OYjMLX2A7FKV3tfhodC2jMcf56HWYlZJDDOTjhkZzjVD3YY
jUNjcqSaLPqYd1jTyZ6pnL5srXNsJX4f53mza2V5SdZTUAX9tLLUlGPCD0nMN13P
hhWx1zvSWhTQVwnN3mhm8n07TqZcD4EM32xtAirRuhqI6awbX/oyTIJVD2tnIfjq
vyYo1Jk843vdtVFf2weRKogmXRiKUah0jdcsobqYgtXw5bcNvJHVda/7LAd3aHEh
HX4ssKxkOqxI1O0epJ+ITeXa5t9NFXZf8P/fXOnL2l/qQMJz4MNekzE/dt43PPJ5
QTmolk1KlplPCaC5HFvyob8sY2bjoyDWiCP6Cd9H9fPd/rYmD/2NjB7OVTRoYaJf
vzYnRMoui8vLDZYLw3zzQNbncHosAtgvJadaTFTuimhB57o9F0lGsfdO7DfXeBIO
uT/aEJItvV9IZ4QWUTh+fhCewatx+jl1g6nXQ+xK5ju/r6L1+R4xtlZrJddEHd0d
euQjhCt2O/w5fYwf7azF6Il8BwtUYAKbQqK2PlHsAFzV5HTgWitJ64+txYc78Pc1
A7DwDgSzMNQXuWYPkqTAlqYm3sKDUFItn4+lCU86URa6ma3f5dPw4UerimQ2SU1A
tsR7V2JdbNV0ZhFnhSoZGpLW+wacsZctU/fUkXxXfZCNTNCx775TrR7C6qbrQ5zq
ufi6ncm9683B7B5EcLbEvKGTLZGoVuguXRCHZZxScQPAiY796iugx6vB7JIvZxrH
wz9Ji8SD+bvItC376YXfppHnW6M6168UWs9Sw5MgK4j4ohLQCwaocv0nX2UJTCi1
LCZ6yA/TwL+wB7FFgmele0r4uoimgJd45uf+L1v7dOKETl0V+pDWqGal67pkSPyJ
fqfCz/E4b57oDccvHSkmLzDAonT2djQz9qZiSZfGzpog0ptTzwKR2X6rZ6WIdRSP
N84ENQ6O2bnb9/XW5jRIt3tRmhZpD6nEJCqkwdR1aN/0KVwU14DrNTPy7X4ARtN8
kOqMAQRKK2biH1ZwJe1MH90jYV77XpyUsXigH/oP9JpXg1Dly7eba3VD6bjMN4+i
GYvwtXfqKVS+HhD3WbKiXbymaCZR8xJmEuE2paiPsz7OPWoUnxLjhN2MGuuvv/3r
hnWHS9KgyqzWSFr1hmEJ0zqbBnVccr4VafSp6vUQOX4/gP0tkCYdDey366kxhTcE
HImF4etXvJlXjHBGXMUuQ/s773hdO0eWGXWQnoqLcfmBv4i5cDRQS8Ugux4KfCuF
pIZBD1ecgWMZjFeXeLFnQfTOetxjRM5jRUpErItRlwZeQFlbxhIFJHlC8n1YWarL
0WyIBSr28sGyrv/UgQmwXWqHXAHfUsleGFhSXbVPdJeRzpapuVF8rFAi1OspTGQR
0dnxVScdg3QMxJAxJinRl/ruo3E1hRhuvCmF4b1wUWB2SABBFxpKbW6cj2IZZ1/g
dKb1WCjKhoZHiqtOqXr7leuenzVDGBSaw3grYMXpFFE6LTa2LrMq9h49NNLXrJBp
Nm7VGIKQKaxhHe8GsNdEKqmTraDcB3UHSAjR0dLY7kU9OjeCtiELbUBvmz0KMdJc
lePO9/SDLFhGijZjwYAZmF4tpr+5oUIKW11pHimQTtXC17k5XK3wiIqvjftu2g9E
o0iCCLpceul5LMP86N63hpDjnmPvKvbHgpfzJOELOovIrnmXxc7sNwofBp7rNqg3
eMcIk9eDomNCu1drnRtyT0QCuU+reX21zNFaKvTWUI6q0SgN68g8cibPR/s6qxxw
KvQ3FKbG1BJReKs5eb2q7eXXGL4eQ3jnLocdqM/fp10Wuco9YwZi14ArWQieVxBo
m1law3wV02DpoMVTCr3pkwR22FIcTi/Awf/5tOkQI7ckGnP4j4YgiQJCTtAOL8Fo
8Jewo6zClMDCMpLdXUS2tQ24EWud/hpfBNSXPQEJij0uXRZFkC4x65B9rccS0XSC
8T0SmjE1LxBSFK7uQCFrb6tFNfevhDO2dH6EqNcvhN6UEafz/ejq9ge07wCn29P4
7RJbr541nSiu44SA1EZsH48jtF/hoacrn2s3xsLBi0Um1/Y5kPukym0ry7zAU7B/
KzXnxWhD31Bd5bg0bXg/ogfWYipkdTzolxQTfbHoiWq+Y822ueg9mKJRIozFFV4m
fZRLOXCxet8UKdAbAqHw74bhBsV4s/1xhbkJKYlbc97PzR82U0yofheqKVC0m1R5
ML3zJHJJdq2pnYIaylLuJ3KhkMsbJC6n5Agaq4ZQyJhJVr/2nuYRwyHQOYPrrzN5
62O6QG96ALO2y0kON8Jft4jYRh23YgQGeYsZhF8o1C+JzvVufJWSqy1JmH7mTnh4
kkaJCvYCtKMr/PzcCbELKvy4NaHoyVFggkL6EwT2QGy+N5bkbQZdhgHCC0IUW2Hg
LCphGA1xBZsxW9b2nvaVmUxUj+xkjhz9byTHKwNawXiXX9LCiY5lU4G16coRzqM7
7eOOcOXeCXezgwiA8U4GBhM0aOhGyb6jjk92QxCp0nDB4zP7AkZz5NTFx74bvNmw
PBvuNOYlIE2YLkkhg+0cbkdQp/41Cgjeh02JBA02OVEr+2gEvH8Hu1Fs8rm6TT7A
QOs78teetecoqOcmlKP93tFkx4GpGSRDOM2XZQAC/U7SsOL1hBbfvdLAEP6XLAvM
2UIHWTdbsu6DA4X3yGO3YYwtc3CD1eTh5SEbQDXfFR4u3Z2O1hSCR4ROtlWNe2pW
kOrBWBhhrp9Ya5vbvXfpYSWLwvjHyxcCE6ADV8WgAt9LL0SClHcvXGygCQK54JkT
ZwmEDyGu0nS9MuL6TY28CXj0qDl0c8KXTiGyLavN2G0GSCex2q1d6HfH0hwANjb0
0XtALIF249udP0EiUfnYZrzHxO9PfgpQ8ydBrp4paEnM8vE6YdWOK5yY8KSH8kWi
xg6pxLZYDq/0Zqwi95aWLwsG2dXjwNtI2FJp6henqAlsIR7gEiWPLrFzTcNXCeU5
CWJ0QGkpY2WihEPF2HudGWEDWGTGjGmvijSsPEdpEj1LJaemqq3k0goYQk754uS9
bm057k/lqbAsURMP8bmXVH7kuaXDO+sRUmYL86GBqoMgZTiIyR6fw4vouflW8vJI
15GtV6vBARyMbmur/8BTJ/D81p8x1FYbQqfCh5mf/HR65J9vUzQ28H8ZchOJPtse
NceDfZ2IdrBm4LkKiuuHnOuBw3v0jOyAyyh9V744GeshoavwCeYOLgaS0jtoOjeP
tAW3eZuOM5SI/JfH/nohuXshVg5sS7cELi6/FFMzb9/fJ4/fhlAZl2f905OERaUT
WJw7jWLdYz4f7XZoLxfOvyfOCKQeWN6R0QsY9EsiRh7w4QTPpkCQQr4BkYoh9gQl
9l8hYimtp1dAyIDEv95hsakXIGKl3PQtsGqEiI0dH4gQXMI6fn6pvtVhxMuhoYie
4dRsMO4Iv2DAjDhvgjLemwJfcV9SBlK8fIXCrz1Oy5LbQDfTTxEFJMwvsc9dPvzi
AIyaUix7xxPi8Tp/oYxQSxRQ+GYFPxnGXoNRuY2+vVen6O6XnDMMhg+onb9djR7E
+2/218U1OrDmaB++ZuuM8r5kxof932OUv2h1QJ5Buct2Ym0oTxqblsrPBjGBVpf7
b/sIGrdfFzr8FbDNgSgdP34zxGD4ska/t63BSpORaqXC7hvSaqnIfL8t6qgNCTR1
JdasurFMnooGBcYYYReuxm9VmeXkl8bpBHQEmYKtd2lQODA3BdymVqaiMOruUSNP
Fcz2wj5j1lFUBvaWA299OyUdOTiorQH25Q0GnYNjVnMPBk4zbDQGSHm6Euq/pGr5
JW4tCfLQYI/wzHwAQ46No3gKtKgAGG05YkrxOamw3Ej7ll1YkclhnvQNlw01wSv2
H34xugR7mpR8ko1D6dFZVUVEETAKl0Y2+qvq8qgVKGCZ+Dw/KK68IcfvS+84+/iv
uenkqd4/Fxhg1gqRwiQBRX5nXgwjMuCPeN+WtwEXxcRCMu9/Thy34WKp967XY76j
DbpolQVXsLmzvsQtDHbvMP3DbQuU68lSzDykzBwmHZ+UOdo7bXlmTMGeYCqJx0Tf
AxlrN8nieaFnfKetsw9ufX4DviYjEtO2oxHB8Xi9sbHk0RE4VORhFZ9QF21YNXUb
jm5QoPdguFDia00dM3X1fDi8NUDvWwCt8Bgj+7J3h2mAqKRdk9KHccvyCERXb1FT
dISvPOXxEDYmcXyDihZcCWfrJhMq3fWzUm9DUN4jkieANVVKhFK7TwxRtekFVqoK
VdRtpJln8XOAgUR5RsDyaAXcmHAXsJ6sz/OrTPjiYDV8t4S2JVgC5aBZZBb2th1h
mDXTh1cG+z63YoAIDWMkEtqv9reZxEk+IlTrg6f1suAlI5icUA8w25KoW0QKDeEI
h3zlWITDU4VB6SMug+KrtdgJLxlF4Zaif6pTowxYBZzxpTFPcg4qOPj3mmg69mb9
ttAu3cSkluF61icoYYi2AeP+o0AF+NMEzMDS+fMgS1mTQTDL81gH4jNkpdBwBp6J
aFExg+u2Ozouq4F9RwF3O0/EjBHCB2ZpsH6+9Nn0WoywcQbzQ64yuVWEueNhas33
bPQx71SIu+JMC/VcK71+Gf0Dnqm5iV4EikuiwPDmOBN17GIlUcAgi6ofvGMlGutl
V24+8qB1wIq8OT34KK3GuxleHb7ctwlDt2gtU3mHh2EswhbyzLu4VKthsANoamQm
9HbUCQ1OlNjLoezEPO83c4jXDZ7RjH/gver2oze7iKkPjKlJGzcHiUe/Wv/Tr11h
fDb3L/N8HvIfDqSQZuTRtwJdh/7pLOlLDF54jyZ5u/XaqWdUG0nA1d83ReBeiEL3
V7JqOAeLQp5DoiCpTBveaAqgcxtD+V1/gtKFAwM4aXFWfsfInkHofi7BTvPftRrt
Ooa0wLbrZgf3IwoAPursRQfqr1WgH5eTiEjG+XPx1EZA9lTxpBByjfGErhwOlnGx
ufnVroGANURqv447ZdNj7JT8AttO/Ub4Kyj7nck5EYoEPI3mdnkNAYXsJnZVabZJ
vLM/mT7C+8io0xHv2Cqg3iqIwOY6PobrQoAPDyZsYTFpqh3yhOnb/K8u6/9A+efZ
YINYhclOkDg6ywiUSxeUJUiqxY3mDdvFF5xiGyDZ6+gdRczr1l0cuM2GjfrtRuLM
Ukb6lJllN1uQVFgh2yNa2JfRyDT0abRHft7RZ8CaaePdhDx5wiLbs7YzCvT9t1GP
FWhdcUJUlWZXRG1EfbUuEw1tnUIeAipOkKN3TDxm3Xpjhj51CvOO9Ijxg0wf1wJ/
IUjFTJZj7zLYMQw9VW0InOwDafDy7gvqHj3ShTeBNXYW9eaWtl0JjwFfL0AHxIq9
sCFDtyf8bKOMfJoaMHEOTGNdQr6mTnKJuS/7hhNXCK7NPdzePkRC6XDZZ6yq93QW
pI1foMNF/rkQDEUck462mZ3gnRbnT0YIY0HcqCcEU0RSj6u8br9OYnLRdLYa4KtC
ZURKRmICIWFK1+doMfGH/qG6cHesRWKtat+pi67yQiGe7cJmrtQ1GQxwJjBFwgsj
Kv3Wr48+RAa1vmsp5m+QKNGI8rX4px8USObcYWCqRks2MKXyzV8HQYJivh9wnd+x
Z3iHzUjfoqjK8l5Yq1txFWOwC35MM9HfxSKdUkMd3vNSgrQ/EyITTloEdg8neUcn
6jjDP+Z8w6fPBedyNhKtpDwpfor0t3e/mIS3RHsg+Kr23AAHi4JAaxBEz7aUssnC
h9RQCayaH8ltporuXLo99WLH5hYhxMZEvm+PleFHijcKLQR3CNaVx4+RserABJzy
AQrYYvkYfP//rWDZFgq4o0XCyLy9wlFAm5PVuWDENzdAweI921J+P9Jt0/udFr1e
SE1ZiZeaifKt9O8KdTBNiPLUaEh7VeOuEh7t+yU4wT6tUdrlEq9FSHLmxxzSKPzO
zQCcP4DvagFSXKa2ThsIFQyEiqZtTHtKks4Vwa/n1sO8buZ5ejlwZxbY7hrLq5yp
kq0yKO9hR8gz+CXW2hBkw74rhQ0xb+p4ujFEd9lWtoY/gcfEgD93ZmvUc+rLw8q2
Ffpka60bWJb/m5sBmzp+8KMJzFlXAl45bDInT6AsCVS1qNg06tCL5JzaWqNaTbJI
4MoVl5Ffp5HkR37x2g37hdnA1e3pQwf4XJt6b1YwYlwKjOGATSg0TWaNZ8W+sTmu
q4+tnN3d/YP0XxzgN1BaWPPO7N70xqftjT9ovVz1DcQZxngePMMaEuN9N3vSN6E8
t3gW4Yg4QGjzU4e4STzP/wQbQmRiIE9SOWgBlmYBZ3ZaFpsBtsguBQrG1OR/9aTv
VM9no88T+/FMeANgFGNpFGB8B6lOkE370//Z6Zv8YP/+B4aWVplJS+y6r09WMj7h
zGaS2gi9EYYAPBqDdcb7qbKcNvM3r+msuQejbVgyvz9bg6JBO7JjOYpxwkECuGlR
fdOtvxQxAMrW1y8QaHp+jXaKkPdlpMyV5AyvSxWSBrJiXDpDiWYwCdU/wdWFDv+D
nZSK0Jwhh7hkYWs5K7RrahXNQqRHTF7FD3h5r7/5ZDb+8Cqu7Ojz4FZxZ+RivCfX
h5who+CMhDhF4bHO/nF5Jw0CP66dVayw8CWYRw/+Nd9tHLp//FZIeDrPTkKSsImF
LeFIa17I07hj87sibRbH2jvnu7IBtq1tTunwygEoeE+A/QFEGAdZs6jgvcJ2FVjg
54cmec+tmXra+iwCdoWqlIB4zE9oiVHpScQXeV+hvw5rDqGdXwC7Qcp2AkSTuKmv
tCaI3v0gy+cEIY1wKJJkqAwCRvDDlWsUsFlsqnwrHIo+LpnDK2x09SnY6Vi9yr8c
otlnzDiG/j/51qkD+6fwv/6cS+ZLEWCsbFdM7kb0hxR9WKHwBUtu136QYMVADIYy
leS8Rrv4cgPQ6N1qM9NAwt1rnp1Y8Hekh68cGvStDwX0B6nQ38micUf2hbWfe6h8
sjhdgGbmKT7ej1HMsZmJC48RpN5zb6QazJbXN6LjnPDjP4azUrzqnvPDXii6qJ+E
VOB4QEWZg6f1iBD5LsJW3U09b75pMU8MHZLqqpd5UbPraPyI6DURSAwcjfb2Azrv
x95AtKczDpw8D8CBUkVmaPFwqgTP0A3B8p5vjtJCKoXgv4xtgBcd41OEzL5SOdyE
hNVIQ3pql+yG+0SOYfaW8i8jFidmu6QuItjBinQitdw0C3ZibFyb0RJMFUKBTojD
2RUyyZPz5QgcbPtk+NUvC3A09IzN5UZr+PPM0MPTXmGU74/EnU5ll7etUJt6mw5y
Ph0+LvCcBEKvSD2AqvdW2j1m9lWLYUFIThxOq0a+Dbe4DLlFypjPfvmyugnRebXm
t3LQnTaAkVlq9xGO+0qtdwXgjIWyW+WJwovj88jgaGYTZJ0kD3m9GMVMX/hzuOUs
Nv3vNzE8ClmLJf6hVaZvb5JH5Xax1Pjexwa5+kEpLQ4zDLcbj3Eeuw+QnH3Tzxl7
r2ZoeaNLXjArAxDPUNhLFefuAF89JewzwzTIHiwDEO6dorIa/LFd4nq/Lgzvr+yg
M1pXD4Fu72lGpJrBp0QcebRsKh8ILW2oOwKNwJ2+H+xGhTHw1oGA0DvWx9pvIvrw
TVxKXk5rJWuKEvKyPHmnbVsUw0gLTa2qwDtqQO82O0nrc+atM7qourGVUX0lVWrE
5lHsfjfQpnbjbBtlw6/dPuN4nFTC3AU1dWzElaP/U4wCn+3ikFNbftlqlGobcEoT
aPsTVdFQEbkMX0XZL8RrNwJabuADRaCo/OgXg6UZD7c4fG2/GA8ndhLSfMk0Bfqs
CmXRhZyinGCPcIxcz5xa/mjVMaBH9HapHu7yLAz09rvWS9DTKXC72lWsRqSgu1Tn
F2t7GmDjuFcU0+ffY2Wv8/44IJ6AXWx9NM0poCIxIRLVuAcfs82qM3DDZ3i+MWYl
K7NdByC2JyLXhkUHvCdAKH8sM+uQeJR7w8CQcyHvcxqaahN6a5wmjUXvVG69b4cy
kjTM02X/XtEr0YL+xAixNJurcm9RhXWY6fYp4PHsc1dVELnxj2Ct8jlp1oB/A+Qk
kWLrsOAe1hmj+CLmWUNHhGAhdl1evyaD4lBsg0vYBnX7lEy8YLf1Yo/mMTcrOJ1N
f9BOKXm/hCNk3n5eVQ1jroCgLbzauUga8gyhkonZbPUiY//V6G2W27K2HCfjrol8
E+3MOIjikwzH6zoSEXqoXCvszk0yMimhC1WcflXgcp704fP23feBuukiBzBq5BWU
abCMXK+DwkteuVprzkNzsLfK9uTHfkL8pHOFbXXk4eMVQck7anViY2+7WZ4/0i8v
MmFqbGyHuN8KsiF5RY3EnN8EVyFmkZauW1EBLXxUdMJ7bEk+eTqx3EgYropieQtW
UhTl9CAyZmFXrlCH9JSkqLhJ8GTavGHRJ48080E2AN2iOZrJ9diqwLHPKuowvQwo
CVtfkhKH2J/0ZlgEORKjobMlg+Az5Rm6bIHtM8a+xFuy2DRViOYuLXtJyBBJCwN2
2Ok8zuDN9fLKenPN3rj0z+MFDDm+cbq1ZCvUxL/mgFiNyvJbT6R4I4R3f0cRppwE
48MTKLqUv0zY3z6HJhRwX8asTAb5ehP2OIZc8AxZLFivhpYEh6nccyrhydgMgmNm
3NG+PX79ioPBecj0BKWovXVAGxHQaZg2ZXg2n/8kxdRGnJ96kql/bJc/svFpAAqa
WOr4elgX5tmpmiaz9F0FApSG/+LNnYThIT6Xu5Oh5UOwJhd+nJl7qJFaaZuGYfNx
yIkELrXtTg/u50e6QMuHVOfFrxvWnQdM2IcyNLwOLTDAyRDRwC9ZZJ+k9KneqLlc
FFGIrrHjNs9I7goFjyRtCGKKXxKx3j24MGKb1MCO3C+AuMOiGffHrnSy7cqv7Yrt
RoS74KOCwq7d5OAhzfQ2+BSUkbecnvEoZON32WkNgQzmQJRZj7ji+i3bolr6Q3aV
C/WbrM7FngtFMQCxCx4PsMGKZKQWK22slnRLj40BH+h87MilbaTadkG79RekHa00
W3VmWeVUQsXLsVR9biomih+3mBWqFm/l0/Tp3ZeIcNq1uOu4JFswWGZ1bYzeS2hg
kDpa+Chj6IPsh40wJ4jQep2xaNZqtb+6G1SDsjCDjDhJipYXxjRMsanVoVNx/GC0
jXWV0xzgzV6xlWocxaWwN83waAvSoZNGfekiv/MdAfj2u8q4TV2b71q4ZcYmQ6G/
4svRmf+y55wBD3cPG1tXPl7CADF/MR8WfExeZ5b9HYcqsh/9Q9pk3Od/jWmoSI9T
JatpGhi4MO832N19iG+Lgdv/bJBd++CjF3hp/R12l1923T5XlevRm1l99r2BkjNE
+ErfVUveej710rb1CpDaj9u/1W34S5hReBgYSlqLwiwRFIIB9DsFOxqYqYMXSx5K
k56OYnB2drPfEcoPEkA0zaPRq5U+qN8sgrp7CXkKlyxIIj4SGBVKeb9/W90yCF06
TzvZnzqONfB1BAPQsbPDujeNW3GnxCbQqTBUHUEjGXkCqqAR0TWWJp0wH9XU3TM7
8znsOEgo0j79ibcCIwwMO3mYUUKHZugXb3WxZUkaqvEHY8iAOSI0R5pXLmZeUk12
3jABXydk7EbXxpGCbNe+mz42vsVJjs/YfXw+7rxs6eKYDqSmWKSd9AVlA7rt8y+T
IgedjVB+Z6vwUu+ePkgnpTyKorHe+zgV+QCw7tYUanyDQ+QTs6tLvWt5BlhFMO1s
+5x7dTMoaMFDrRp9HwZ8zkafBY4+KbH4HwTLHcg/AYaWGhE/roUf5UnFO423qWTX
Z30JZLbx8YGIC5K7g+uZYypqsVeKcr8cZDtDQ9nFtopULlUQAlBhiDL4cJE8Nvj0
BegPPSv2iborDsmaClS+J6F0i2xMslziL7UteO59av4lLIxSrZfKyv5lV9AwoZze
9sT+0K4bmuON9RRDlmLpXrK43lWepsBEwoG/gW2U+MF7iUqNo0fnUGbYtt2cSwMv
NKPesiafGV0EahvdDcFvjmZuDGfSz6YEDoTk0kKQV3DnmdDRbuUWkOVo0NmES2gR
uEkOPsfzuwlkfeGeynjAag63nmQzdyBsSdQm7UFuLLwCmDPuwFh+0ew/276/T9qV
S4tjAYV+VQ46OWN8lEAHNIeoV6ee51OTsXuB57fSwV2pRW1QGWkUB1eiGaZsS9Rx
TML12D848kBOwgpwZ5JgAeZwa98f5V3acKGtGdf7a+2ntumyEYeDJh30g9ycyMCT
erwuYVE9nozLILvvjAz3X+1AMeYECZFNbQq3Spv3h1PT0N39GqlREDSkQdN/hFfk
f/EVHWx+LJF3FDG+zFQaO+KX21kTihez6wX2F6GIai4qE7dpecNxAdYmYiwbbR3O
zhJpI7k6Kv3zyrPARH0mW8+UADD3H817/0oIoHGitCCRcS1PC/To1b1yfF05AHKp
tpqD7w4qijB6w3ER0mGPor+Lhd5tD1tUmNMMzrIa6gsFkoCMLbPd/km/trFt0Tvd
5gyf9y7G049xcchfzjRlYz3d5PjtZRpWeWf/DU6Ad6P3QW6B37FQoNR992jua5Cb
JbPq3nm43MKugaQkeylEszJu2wgmH4sHYh2TluV+KCTsTU5CLtJWr+ZT+/HrIqIt
qkuCx5Qc6TNK83nhYaufnKyaNTTFNSbwf4tR1CCkdmueqMMfDmDeRqfVPpVOHfXb
wBADF8CDljh143wGPzIjr+CWyunyD5Jv/x4xuf3BoCy7QJt/u8nqiEVt8CW+0SWk
xSOMYQS+Q6qQAGjhB9vetVKLWP4FqhrkWgbhId/xiha42lrtfK1J8lXHXLq6f4xJ
HhlphLHavF99fZGP074R0J20vI+DouU1efL8p2ZWp5UXQJPOsawnN9qx+hO5CewN
YH42FGq5pEpAQ4ugGVC8wPt0L3RcVQTa9JPqgl9tmDNkH/3xqVAWiuGoudB8CQEz
BnbvPo3/jPmXvGGgtiOgb3srGevdNsJJWHQB6Me4asWVuUD80gZzBFPrPf1hyg/k
ivaXngK7TKRZIWpf+DkVhgaKQlxbzbgoMQxD41gBvAdLt3i8/AiYqA3lqYOIE4uv
UTMF10HVsn6jfjE3Xf/Xqc+tCmYKgdIpBvaXaPcbP51FV1H8tV1Oc01XlWjEH/0x
iL0LajISpwMdt5ClCqi8oYwcpm+SzxJWgGptkr3oHsDy45XLXk5hEXmXhcDahZIr
/JBvu6I9ZJBARstgReyj/T1mncv6c3H3IYfDaW8NIWj4laDmj4GMJTQefnFl73dQ
2up9UX7S0Dic/sci9rXJXjqAVi+CDAAoQQoWuC6YaE755f/8kG/lKWBjhNtmwRkz
lc+qcRspu6DBKuiejefGuVg8z0ttApltifR2+Gx8sTXqFqXn2e6KFV1AVTie/sEm
tXiXQRNAM25WGXgLS+EnjXStvptqR0UmSkyeUnNeytma8eoE5B3rlV9PL2kwvhSA
AfM4QPoBcLU1WMKspU8h/sONzm78wXvPjEFCA6S/uj96e0gMxJS4Ko+2hJcJ9FU0
iu86IrwZtNvVG9Cl/5vwfXOioGztOrlfLcpZri977B2PC0zqvNvYVrWUk6+OgF9w
DaqU5iKSK6s+RazG54AdFv2LFFB5BnRlIHiKUkcjnMLLQ6TvMvpwT5vzY99p3oaQ
3ptZIZq9S7DNdUS76uUydrR1M3ubyf8wwBYhhNm2OaEu3s2BEDyCZoHTPp0vcXue
PV/Bza6n65AOBL9y888cdhmjaY/h7n50LgqnUZc3B5Nsq4fI0xMwxZvaU2vTXM/k
3UNXZt38jJD/TJPJSHO55rljRFDITL18HFm5625SjDLw53IRn/hsEfpy5RkkjBpQ
ntxb0xmfm9VbW/c9yHBde4v37YTZa7FSy4hZVfiVIkP4ajVzAbDp7S2I8T9tHDG/
m+fOxOMCduMZR0+6B6g6m338GyykknaxeCO16dmsCDvyHUIegLdUIKbFATBZLTZ8
s83bKBu+KN9I2Rqo2dbLTkYB61ipffYdM/Arwe5GQdQEucZALGj9CIoYFcNIUgsy
ELEg0622Cmn7qn2Lf3Vrq3/20Do66BE1F0cHMkmQllqgWH8pT0RYcKcNUcbpRYlQ
C4H2Rlk/iITEv6+JbokGGyLAHo1K9c6Hok0X9zZogDq+88Yxl2/3iJEQHPT47Vv+
vcBJUOqJqMtgLCFCF4O9f/HFHyrJOhfGuFrCcACsuAr2l4Ebd9GkXtN6ziqJsV89
xpfG2yV8KV7Uufe2qmYQUNcOWha7XvX5i9NM0L7SGZhVr4HRaatryTCYTV6kkRxN
DsJhX8u1RUW8cQm6fUstLV0W4A+H6rRgf0rC0b8FMB/44CwdePic24W/WBIcyYkd
he9dDZUBdocULNGyTQVEFcfxpZBA73q3B5Jh4285pwAQzUQHCP4WXiWxHkvM6Af6
0vj8yrjhyzPXS8Q63Yd0O5r4CVJJ61mStACC6iR/fEzYGLL3884+xCi9utweh0GL
N+mUokllZXzYW+JfwT+UIrxb7RlRfIvCCtUO7EbBO/JeyDIanN+YEfJFoNzRk6AR
5Ok0d2aoN/xcLTpOXKfWDD9lazR+eZ0hVu5LyXCWivEx2rzBbPITqe+DiZebEJD+
5NimkfA3VZdAywDPjmC+eUBpQ6ATJJm5KQX0CBZD7ZIt7d7qqmdWWNkHKM4zEe9x
Xn6qzTBIBhZBRT7Sju9iEa6jRWT17RrUgd+hIpmSbsxlF7gISJiFv0W5RA9RS1lZ
R9j0cWDsQ0bEvNXcA3/pOpZgmhbsQ7qthzY0h3GyX+QlpIxrWfz6WmXts1FOPtlF
JIrLPVZsh9YWHkOSgr0s4kQaS61uq86yc78pGP1rNhyZgjBKGeMwaJQBY0jTkDNe
HwCGKneNdlmykbIuiBQWvpMekN8Qs1JG9R/4s8X17BrcHFvzgM6I7e+po8qMbeiS
H1VB3AOwJ7sUhyhs3UMijCGXl+tlV/KE/dKOKInbQT3XOsnRQWG1SoJ3GsHu+JCg
Av8oAS83Minpb3csHEL5sFPyrIFvWf+BXw2+rP5z3xWGgl5t1jv6fB4wRn2sEv9T
pJN5Vv7kxuEVZVo5p0ErUXHrV3e80SOYBesRp3FY+jM11rcJKeerBHNoRtjB7Ovy
q5GDhzTKZiSJhIPh6jJPZKn14F85r7Wlvwvxf7MP7BzmNgUWea7qFhyStgwX2NrH
foLNYZTF8cInNUS9R1E95WEiugA373GFUO5fd3iM58HgwuKjFd93+o0REHJcgpza
D+EoBu3ar+klaHTTGI0rp1X5z0NiJvbX9lz0Q4xHE2fEGTHbYE8aOAHv6oYhWWtt
/Ys76wLLuOq2qU0edZFUAGQ7wP8zsvZRK9YEtEs3buRhr5RF73ni0SjXnVHhJiAW
y0e0F2ZqWd+ZL4wz6lucbW3UmffompnPbqEJI++3GcIKJ6waJs5yZ0A9hrW7Epd8
8Q7wMIFXbCgHvnUju3h0O9AO89krsoriwYOpVsHLdjYuXFeziW3n8n7nPf7VqncJ
uop0DGBMGNx+vATbfK4VNpxgC7aC6HSeOOnSEYBThz83E0dHuymgHAdvvM/clgAb
fVWeUONustbb8PqUgdJlIKb77XBwzhPw6R9SyYZH6S31H2A0zWpD6W/AVq/Ri0Ib
nFJSm0DtWH/vgqpXb6lpMkMpzTZnEQnXzgW7ZgGxDcQC90XohUjz1LAMpqWtkxdo
8s7u5ifG/xut5w2BoprEDl6yJ60D+2feRuAKaPHjlfEVZ11vW6qKCgmR1yzXiNsd
I04ANTU4ryKOE1E/WX+ICpaur+6As+6n49ObrgYV74sI4+TUHo9BJlgrCHdduTbu
dYLUs3z2RCbOFQzdG7UaqqHo26E6vXazeGoi+rhJyENDokB7GQHzbldmY5ezK1NQ
0ZauTYTJG8ol/ONPGKPM0pLdHAnRmV5isewQI7+3aegnOsVQqICeSzhoAqVZLfs2
41Lixxpxp907LV+4MDDF2K53tatbv2hMhqf7uKkDd8L0u/EU8Y45y6ePzvs2u+YY
OrqjbpuoCiUlEHHffb42epToUavNDTGEG/cPTAhoWObWpXM6QRUsgnzWhgq5CSLH
eLrQO1mAiVnooBOzxwRg9i1eFK9UoyFhREGHu3z5wSU9l81Sg5X+5OHs94IQp36r
870cyuBv6w8w8gMy9AVJJW+5E/ZBtCDA4Dd43DUxWYBiqTX1pdL19zP8rTG/eAtF
Y0SUMAZqH4znLg+uQP+Fhg+T7CsKh0MyLsou8aLtFq2eSbsDjs9Us9R3dJnpJX63
erIuigJD4106j0Oxx7wbDfDEmy8be0JCLPW6TbwgTJJiF4TKtFoG4LFdNU83S9mx
PrOHggg+iz+g0PiQr5IHqDhsiIAUg/NDhsMKAl95d0ROUIxFxHYc4/B5+s5Iwy4n
oHFFYa/JZ3Nyj45i047ibclpf6UjfsuDuW5XSjnxNV8g37AdFt6xNFmhzObOeooI
rn6iASGA2q8oiV2X/V1toCiJNztByoz1xEPpoQklSlBYxDW0+jxb05+DtEgfGZBE
hgG65IcmlIypqHO3jzsMOcGW6ycQNEbnwU1JeurHrZmn0TudpFEELBJXsgUysZvu
HUp4fInM1a8w5XNqKfE8bT488iAHdMqf65UFjg3cJ+9BdppJVmRaH/xCJdKCuWGI
HC+lId7/jH6S/IZ62clR+Ejt8ETZ1QyP6Pta/fSDnWwMYZRiy7OztHXoXSZhakbE
mt2z6SetBr4Eym6sKvsXhV8X9B6RpO9rh0el6FKpSaXCeiIiqNvFZsjTVvPNrmmE
oAaxMc1x5T7miLwZEVDJyeEkSbl71CmePVjFflXro9DgMfkdwRKYwX5BrDaC2nO+
m8GueZnhtjGPHpzvxT1xOe8VzoKmyow6YjQ+7G1jGNW8Nx7XICWahPrjuagyDJF9
97NSCE80weFqbEnORZbJDgmzrPCjHefJmoQTuvqgCR18rLa1OFTmDM6yH3vNOw7r
NVmT7HGoPzEQw7WqfOubcvwCYpJ3wVaHrmq+3+h/HcJJmJ19AhWZm7UpjyTfoqwK
gbBfIG8uLwxJuZoZh8l029E6aNVKplx5rvT58bZhJ4eYzGKPCdIf3GBAO/ZJBMIW
+j6n5iWGTYL6No2q6DXFqlHeJbK3ACZx/shOQnpRgCgbYg6c1oeL+la+qvl56wTM
0H4XLNTdYJXBF9OPHqFyULyXdLBjAMnXMyoNoTJCDohFnLi9UP0LSUSxNBmqSU7J
eBVzG/C7pHDdp0+Rr+hFGXcNkZr/QZiHj12uqDujhtAcMMVRaanbwZ12yYpNU26M
t56wolNTFVq0Yrp0F3arWiA5HbKfJdP6vLqVCkN1VEpThttdhg9zqp1QANIsZpVk
ImSZlYF6GldkDchZw9RjYBtMx8zOivB8+QcJBfPRn2btRnlDfz3LN5SSbEau+2iM
wFgi2jFDz+zaz9ynPNjWnIW1vSKgfuZNsEiyzMzDV2qJsk+KgMR6KbDve7pgozSw
X9ZLowxDHsTKkj+GBzpMhy/wZ5rSTEVcy+F9hd8oHS+Sk+NACxb8AxlIuMCIwl7n
hwZJnDzN4QGVNH8IOphQohUn86M+tBgfnvU3Da3Smm3Vywi+lGtGKF/TiRSQbICl
mkPDKt4hBjjpKHwq832QxdzIhIRp6wv400Zh1avF/80jE/VON2BtiLFJu6IlFAcv
oaZ165jeRAtnOTGfN2JDgSyzZ+IvrAZVfgQe5Ub2+WNFvoUv+P1n2grc+s8Z+Zc3
WNElbBf6f+J/ciFUATFfPDYLNhEK+9ooLfi+ois/0086VsMPrJSWe4XaRUEeDciO
KpcKtPeMJ6hPDenEvssy5LT9Cch1pATyVYWGD1DDP+UAI/S9REU8FnJUMLa4L/Ak
CwKcXGzliCeM53hVZ6bfpgpVLe2JXoJ4xD6B4+qx/2/iTj5T/7LGhMJXJz0h5hWE
0+3L7CkYIeXqcoMQniNbr6FzK4+F5vAd2NYHqL1znIbB4jRcJ2mzXTKbSH2v9U5X
60+fKTUGRQw7MbBQIa0DmFnhtMihNqE095nY8sinhmwtKIfgWE01CMWy289KeoXg
BC7qnbyv0SHnHSkYTL5vnZDog82ZhdNXMrcZnpsvuZOX3C8tY2NXCmGOT8yZHYvc
3vfXOAxZp36j3GWAw7fkGzGcWX0IQ8f9HDpFmMoLW7AxG1CEqyNxTPsqwppzZEAy
xOQ1lAWAt0DqgAcnyXXpbAcP/kxdqb22/Nc+7BhvicmNU8+OBJ7fwS7Lp/Au7odb
pjBEXwF04tuuK8E9GV8XwHhJP0z80LNzkgLEG22xzLhgKHDSBNQ3MNkjIL89TBUR
dAM000ss27JRe/KbIfrY0UykA+FbA0xUnltKuNVlEseD6/bTg0LhWJephoj6tF0U
icfsq/+V9qgO8vosQB3A9zh3GYr5D5DegquWHYu8US76MTAgU0i09CEDRSl2Rl/3
GdgETfgiyllhJJIwqnBIbXVgjATa0vfBQScwBsRi6ZHhnUIKaVx9cERNCXimf1d8
pTgBVykCB7FEYzejhj5/99PoIWp2X3+F8Jp23vuPRx8Wo2UxELOl7VTaLeaQpLRM
biEAB75jdusQ+z9ugZEMIvd+wah+LltxUAMXD7i2cPmgTL2lVefyEm2gNEJaNYAm
tYhift5KyMucdXh1m5qkTkhZMCpNoE44uzEc6yvlV6+vEQ/S7yPg2qHjA6jP5Cc5
xypSiaPYp4BrbqbFFm9vCyI7ckaPAxtYqNzs2OCCR2QZJfSteXZyq2lPXcjB6ysF
VS0GiAkthlOZ6U8HU1RxN4iIs1QTx8ocMBHJCAa/Aes/exGbLyKPIne2X03/ACOL
vylpBDxi8zlg/RmQs1pcbBHqRBWl7E2jrDdqiPd5/QBprjl1nX8B509LIZa+UrxF
zouaSG1PQk0nRWdkRwUreEK3t7o2eaMECElVgXexo/ZlK7x2hg39zpBEBaumRy0P
mM29uebquazB3I3AJN7uuIQ060/e9hi00g2HxVtVUMhjh+nfWce2ykqUxCPH8a1p
n5wy6y7Q8Nd5E9Of2NI0h6zDN7upZ6DBwc8BEjWk+cBuiOig+aKg5rfixJ9LAhxy
HoaITpK8T4Ld6xHE3CsHX4+yOH8lHrqh3EiySZd1/n6oRgmx1CCaF80eLXJoJelu
n1KaXqOOkqaTZYURHbyIksqPt+oLRAv3TFyon5ec/Jt6QtWOVSKReB2UKtDABtbn
25y5MapLK0opHlK7Fu4fYh/xApf81lbCKtrYn+Uc8iDP2rtFip2RKAIg6sgHh4Tj
itMI/9IuL8fCckZVABtfZGtcGN2jb3H9oSf/DlkfjfagBv9vNPBmsvaU2oSUZINI
+/SAY3Qgcl9M9VxB5Q/FgCvfdrNfxVdHYEnM5yODvvgGyIp3dbrbA3CppFmD5Cer
123GfWy4LFwuhqe4s76U8A/pCo9UJ3/ofPCxRFp85cqFA2J93hTuXJQ8dgrguPHH
sHCMB68VO1XJ8OGIFMM+y7MlwOjMIVomNdDlgw0L8LSmETubDCt5lDc3nAVVY3mu
x4MPoR572r1GQfcZIj3MMV0eGp0tgwKWe5X7p4L6I3KlRYWp8jYiiaks7a1XcMb4
gIPxUyaHW95U0gju+T8T4l8sKcfw8B1+6xtWt1m+eB4uLBqERT8oFX4w+nec73Xf
6osG25IIGdsIWuTx3cjEORX6rHBHEtotgXkWlMkNsWynnHKm79dZN5/QuebivHEP
BIgKnWWqmhwaehGx2AkBmz1xCjRmyD4lm3xrJlO/oxhS/V17c6IpFDlOQAVAhZJC
/mS5yUcO5lnUBi4JsTm6BGE3k+XO88YgyKH4OLvR+SIL9H/wZEBc3cBPKe548cWD
m992KjdplM6gICuO4vxrNEJ1LNQgN3uQ41RHhvpcvWZ0M/WLsMHVKC/vlAWJ4zi9
rqZsE6VvZLUGHQ4gnhv1s7nYXXK2uRyYLUPQRydZ/zdAHNwYTUwxaeyYWjae7ADi
OWQ/FyeQ4jh463jcZSIgXOnQJQzMyrzfQzpthP+3mUbXsInfj4UU6VcyUeQ5Dix/
7Sbd5hkvH1kIJCccvpnADgmOu+Q7rBPIIqG+eA/i5Jr16Z1eiwnUvRX9b0tNgqjP
1MudVmxioLO1kdmwdfOYQDVK9DmCP5g54g8MZpC6H24VqsDp7zhaw/sThQOdpGuT
g2IJ2L/8oz1gQpM6FpXvYHjeNRGpUgW8fxTnoW0pfUfGyUxhXEXb1etAMgkwkXYY
qqzOUdl8GAENkw0yC6IBUirRZY2fx8XVzbmPz65WSqimu5J9dZysBV2hO2c19mYr
yYvZoKgp6wB5i84gD3y0fpaEBIDU9IKJua5lpnhJTtnVMEkuDggP+iXD4QfP9sKC
YZHo5NbECCn39i4ZWzSZhqYtiwJgyHAJ8wT7W6HybGsBexU513yPkVrAYAdQPnCK
d7zvy+CtukMb+p/a9nzshELK8A0Fi9v/0nnyjEFo7M2CRexwtv0pvebPj0i47Wu5
Nw9YjUYGrKHK0hd/ze7c2mygYuz3mzOzAERNGq6IHtRxgr7dyAV0/u4EW/ovNQ5d
TK21YW/wRely1LtmQO/CN873SSpIF6UfKOy1vgqxV/2tw13PbUD/HgjJBNy8MKic
Rrt/zwHgj8DmuvbLBQgn8xIgdiKZjqArpCsoke3OHDfQu0ju+ZVfRBvNzLYG/pW3
Pe0jVQn7lfcCsBtRLNGnd0o7arZ54x2ALKHmJ9C4r9RUZtYY6f7LHAGZ2e+bIXjN
0ZrcZVxWhp88RDfAw5/3zzPPFDrBon3iuOAfEljSF68gtWwgc3dplX/OGc9O2chk
9ndeRLIk+yng/qUwn2W1Ha8EveWWOfLRbo6YlGYIMD+2lBCBdrK1UYJihY7hqyMo
dI/LSsuN9UAFdGFXR++93eCa1dkP5H4dEKFHwE6y/ZO7aWJ1XsLU6Wpyhs9c/8wC
BheIaARznLr3Kmx9y47BoSyGDragEV94ZXHIPjxliLhMIwcHk680l9Bt1f2LoT7R
ShJvcMY20b2h5Ovz5dtI+4rwEteemorq04i7oLR3gUdVoC97B8F2rJNzm1smDFu8
zwXcxQD5tkyyLk/6365mMzrMmuWNe4eQEYZVAO5uAtNhsV7jfBUeBRBmDQyupjo4
naWVWYhU7LC/TxTZ+fycdmW8pDevehOR+pDPHbl9AW4aEZANItT68YpLEdvLsJOt
uyif0RaK4TikUo9wO3dvGcYC22qYiSEZyra1n4fZP+hLVPVmmdKJT3d+mcFqFM33
htbmJK0OlwJ4te7N3+nMMmzwqtIeF/bWOLuev+rBF6MkWkOS+MBZl7ZQH62m2ooA
aHHu5732ExxfCXOYhRfgrIhAAQ+hI+osVwb89i2wmRMruQUh09FuTDPyoaBavS5w
+A47FDPGNc1SusZ9QiYLOydKfgH5lFaRF0fABNXJazHFZscKEHcQjBErdmIUwDaR
Fn+bJz7Izgu0ITjEO2Qsy4kUmnsMTW8CiN8fWz6oOIp4PgPkOUHru7zqOdffp40v
IaNc7c3zFlDEHixagpv+J0O1Uif73GTs3KoxqGUX7+NF3A6mqLTFbxzlXwYOpQSk
abdlhyht7jZU5mn6/cUh5WbcLq1mcMkZB+o8q0MK4JhIH9KbaoLsfLoLeRUFgb/c
aGxcExDkg3Ioesv2WWzd8OulSssBNo3zjve3KbcKituWUqJIa3qfhOh/qyA2w4qY
cmfBUL/i8BC/CSIb/+pCTP1DVpuVNcvf3UVwaH8lhG6xYafh3ttESZ1kOdS8fzDH
J7EfGedodNqhz0INSec2P23l6vthJFhJubXBo5UynvEvVRsJIP7hG4HkaaNyBOql
Yiadc1P2zMcUOyufSyw6O9lETlG5A9t+3huwaPt/LCsZ7o6Kd2i928dc6HrN9uJf
cwgPQQrKhtUNaXYExfW6QOZ078gtOH7tMn/IQdezl+SaZ7Hr1YKKu+epDBSgoSkc
RNeR+h74fOY22tLv6xvJMtp93U+L9dNDI5Bs1joc1UHP+LedAlV2OwAHhg17H12k
UNmjj3cfzFR8xcScuHq79aPex0jCD8CxF2YhFfawYz3PQqCFOX0X0HMvvl0DyG85
4mBWMRQi3Mui510RnGw+RwshnX6maM5jMIcRsfFiewde72YmED484grwmqF6r1m4
e8e7KNjgM8o9uzRNek1vSVQZ4gX0ukRRRexnMi2BzHmjoh0W3pqZI4WyfZdee745
Ui25ak0/ClQBVAsJyTwbh7HDBtm0MFwyawSCvoC4OwC96giutwgKmSZsyazuN60H
PSzJanKUOyZc2P0EkXs9+2mtncfoNXGsNFYy2XlMIW02LBFzs9iKMl46JpBTXlLo
5q7B42I79hjQSxGc/jk1Pe5JU7GOXqfX8qZsCJNuckEEqbwQZk6JNraMWFrXSA80
KMETC8LRTeqhCMpEjzQsXnl0DPEuoYZ5agzsfHAysEYMni0QjFsxxEwt6nTYyr+h
8gRGuXSnRAGUpLuaBPnoLGnnJRLwH87xVhtLJxHoq3qf2hKWLoKziyShgVhXmvrK
hhs8o//3WpEAICYFCH6lc84fnUvrNs/p1K/pOjV1AKhyWjNZjrIA437Um3i/Xial
oyAxDFSye5uSgla+HxC+E5Kf0CeZoXEAbSwr9qXvgpPmA/EaGPgeckQJ2Cr7rk0u
itLdDxzZSvPZHJWU4bXO0ZxL+hwSYHnPpcKDy6x39Q76C4WE3ZoaUgljSbqZm+OR
M22hea6nMLYwHACyQssCzxfNoz2wbhWLYnX/Cl42zwklY6Eo67Gs7XCMK9I64tC+
EQn4h1LnyaRpw2zOZ4ogJ0TkvgPJ0VD9qY5GemyH9fbCnV+Kbr+Hlt/aGx8eOf9R
qC46AAv/rc6Bsyi6ngwniuLXMIvbpW8Zx9dQ/SlILjcEBF7DFKd3QVqa5lYi2dZ9
15U85EXS3Vn3jMuqnsH/h9K038sFUnNhsdUO8vyIiFmQbXDn4Q2kbDjXf1atgMAM
32QsN3XzVwkNskE15Kmvcki0dsPXnvFHUI4sQTT/t4snQ1a3UdZh0UflNhlDdI5E
J70tAVqhf+MLxVIrczt3Beoayv5nuYJCE33IlijTTRxWlKwZ4OtixIb/eh7YbH22
cpJld2+Z3qQtZVNCR9ZNKhn2E87P+Jx44X0ZtBKoS5K3PPhs2sw/7W9NaWmbo2g6
lX2bXHbbsSwVjUTWUpHN0DG3K0pON/napnKZbdz8Grc3yFmd752JGB+x5uNDIHan
HWLnGOMo5t3bnqxKjIHmw+eyVDbxYRD/mBq2lXR9n+7f2akYl6MZccfF0Cwqzmax
FVEPmY3YVLFsTd4AQy6YjimSIObZoIkUPNCo3Y6u5oduvgHlWEG8ujeJYxtYt5TD
kJ8NqTAZ6MV/+9IiPGzsA+9Io88b8Pjlmf7PGGm6jxy8uZu99+vzdxCN0s6ZretW
32BXP+QvgmedhZjmE5uvpBp80k4WGlGAILwVq880R6Q62TBLsjHDBo+a8A40KyeP
17ZECPfDDJA+okOJI47gdACoZfDNXlvaL+Tfr/Z4nSkICe4JQ0faFtSzVRSW4nGL
azP3SRHJY5Wl2JRoiiO7LzTcUEFdXE+uKLDNQgFSdM3Qo1VoFhyj7tuAtE6cBgwF
cnQlrKlS+7mdZpMf87mWpyThuVb17Pq6cZxcp2dFSRiR9LG14YKTc+pmJyrSuOPr
VG2tvKkh0Q+stgOjcZzPexOqkpi9YcWgFGjKaZTVr6gBhieDvXg24bsGyucoOTij
BKd5qYkMgV3jqBtq4lTIg7b9Qzj0n4+x9T6IO9vSKPg0ofZSO2bT0rWxDMf++W9p
tN1PTeLz8gtYoSuP6cuoeYAvA4b0zYUV1mgieN+coSo2opvV6Kveg2+evATXNgOX
T/KL9T0+XoxrFptuIFydvB+mwxRBRsy+9alA4wKIwzP9jZjjS/yLnCrNjY8nTSFC
7cSNqSHa4VKhY6OO7Be88dSX2sugqv148KstJmZKaqJfyWAl0XHh0BuY9Gi17UTH
pcpRogsvsNHXs97RcgfH8dyB2+8zxs5gdhuDvKpRmYNWeNGBO54KVRuaIXc5olOC
jXJ/Lrl84ib0LwNVoam/rIJiyPJQYW6SvG+2Z+t8BoJ3A0oEjRNw4sps7MrIozUo
mEwuTyECMFxI/yoOnC4BTaiw3/1DRuk+MKMy3epyDswE4DyKwJJZGYgOmwv+j9FH
M6ug0odTh/5qOuBDbqKkIsBb2DSGiQuRek/ht7vXN0FTx3jLAy+xW/7X3vjcWC57
6R5GGdz+DbFFaDcnsOnATzoh3rEp6VR1KYEY30FhE9LVeTrQe2bQvE74by4ZGf4M
6JSOL7R7VgcqpoEtsKZwyRWaDUskEx5s2xa68stY8MOyozjjl8fSJ3PfT2+p+zPB
pMUqXXA3zuhsysBnrrJCtBj1r9vpzSYzSscUCgF8TqsM2bgYyHrCWehunVcyuEFr
ketJySgSSauCiatwyq62BtkBb7Gnr/8sJdqN6ks9pDtAg4PZydbMxn9hT9xB83IV
zPTLn57syI59nztUQtZul7fWkcfF/4zgArlnSGigexbpnrTABy0+t4S80wk32Rg7
vHtugiIWje0bmxOxpjxb/0oE5gNsw7EHRg140+E5Kb/H/pDi8bWqdZrxBxPCXSub
Hco39tOrvUHsBZXgWOy6gYBFPZA6j8rRkmw8KGJk0UMB3pvCwjiuC+pmsJ0PW45J
ooabfcWjoDw4Xr2n/wDTgA04rvf9rZqrI0V7lN+P6z0eMs4UdBC823FrN3vC3JdV
2vrEl146sQ6uBGJOOB4Ck5ONTGLqjdS8j6d0niHXovLpsulxolrnsuAoY6cOQ/hh
DW9rAxphWe8GAxZozhKbVcFF0/fvxYmpDCV3a9sjV2+uY9mRCDVs5ShWBT0YAqUo
9NSErx/DLvtORfT6E8caG3n2RkqkjpHIFlqMM1QRNJLV/RopMBOx+rl5LpUe1y/U
N8NtYGABmULed6KD8D00lCvWazQ4Qjex4OWUTAemzBZYaLdbPpKEp/ylMCNx6BYX
OWSIJJMx1fV7GRUlWkYtdSaqZRhqGsjPa1iTCwvy0mVDRiOFDPcBZuLpT6OpqxFU
vRoM7nFJUxRM2USufp3XJj4UzOL0yaL1GO0N0rqw6IZBgUFyBMZlwGmGnwNFH2+Q
rpyGEhpDm3ncUwLs/TPunr2mkimZq6BXIx7vrk/k5UI8Gb/NRegO4Co0kwbEfLvX
ewdpvYtl/+6JnktrFAhi3cILrcTBcuD8xqBI09JmBkO6+ISXT+Oc0UwjEMt1KCJr
0402Hj95utQyksb9BYNNDe041a/w5YZy7F8UJmA/LpgudyY8YCxDnVKKxUSp5jMH
/xVU9jobU9E4RCX952KTQfDnma+Ehm9ky1yW3JHdujXxO0QZtiL28LtHZIaBw0/z
tY+HLKg67DFtmT9hqeHesq3KVhp+bmal8/vl1HBcD0h79GFka/0QoJRjOtS0/olR
VpJcCq+KYThs9fiBY4Hy3kqNKP31CqgdJuRfEGNnFB1OuWkYCJKrC+1WURPVrL/P
gXzxFHA+NTYBqP4OP8a1IeOlja4vC1SX9VPhexxjD4GGYQ7ahxYc4y4SokPb0qEC
dKmiaVloH7cSOjJwmjp39DG9iCIB2Q0Z9PK8HwJ1QafKSCN9+DnBIe/ES5ZxXIru
tzq28svE/zjv8E0dXNIH65hhOC8FYN4XrIeQgcwvPcjf6z6IvWACnF2NKOPkNwZx
oHSziApbqfiHpn1NtkHfwa8y+c+rgS0l4pt9I3wuQ/kjebTQw0MxPJiIp9OtUMqZ
HS0CBOdBp8JW1pct5x3jBGvBwrG4nKtFUFSfs5MXLQp2F7boI66WBwAZjrpdRQFq
vCM5QzGnPiie7+jyNlE7XD+0L8WMsLAhHM95WrfZw0DGqpAvl9qoir+ybKFR5myp
PAj79QfHkPmZTwd3ZT7LEgKAbYMIgfIOmvy6v6u5g0tKwR/F5XyV+PX8XwMU/ZfF
BuuHO9atAxpB7Ola2RZRLZm4b/ENNkiNJIAw0xYWp35AISB6rmnO7W65UCWmuizn
qsPgKXWnbImQP3R1W1TCh3cMBcXnlfwxpM4nAbvBuyZcJ4teJtyK6QrH4XIi+Qyh
Ks5mRzSxvfOATsD5zcLMocvDfYczXyrUuC1sXKAZhwyk5Ddu8lPz1lX0ECbHDhMw
yBgRiPgk67nGeksIShfPmG6xZQ9y/cmcDSPeLwUgzKxXos13F/lREvitPpFt5PZ1
T914OuHa6mWZwJjDb1og7ElOEp+Xo4Vm123WCnb0rMn+uDXtm4TLFAGzic6p0znJ
v0cIAkfIPyN1o00TPkLzpvbJFZmR2qR89Le/+/gVFuExd+eXf3FeTdj6Cwjml+oI
M9cwCmBRndkMG/bdfNwiiUEr9mHI4bLT7pOHIAkflZNw/o/ff2s5YVLJLhdGXzNG
iE6jZbhUpeazu8Sw4lIGqCEcCj9C75KEsZooEYYZCYSJRe5Xunz36KEF9CIBLM2b
urpFQTfVV07XiQJhZQMx9ACoDSdv5ozZYlGeiiPXQaNj+qT/BX6YtKvy7nbkSesS
Bomw9kVvsRCiTihW5iEyU5vJpd2RI/880p2lItUIM01SqnAWc8dw74DfeCw82+xX
Wj8o57ssifnoNPKWbzPpv+DdG7mO3enktdoqj1jJnE1S2Kh7fgN4kvZBrNUwAp74
SsXRa+US3nNh+b1oE5i3iCHtJSMlBH/y1vXWx2AF+8IJR1k2uL9Zr++SEXNftj3b
3PdK1oyW5+LTqpkqN5KBMsg7jjIDfLG/CjjMvVzR9l45suTYQ3FGWCSyL39BTIcs
NRV+dppra1xmkfGVBI/0LU4d0BajlV8z1vEkqHK+G2A1/2AOUdZE0qdkHPdymGRw
cRfZn8qv/zUpda2EABKBiTCU1mOFpvX3g3kK3BhE5v/RFaxW/gjwZtpJVKVYlMQP
`pragma protect end_protected
