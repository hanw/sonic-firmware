// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pZ76AM4EP2E+Z6mOSi71ZFE0RvttPwG5tRQMZm6we0RN7+BDvnD+7ch44jSHUPzg
CWpMcXZwa/RAjjtiq/KaKQtNrd89MBHbM8XTAtkZ5RrVgpFYtaweJvXuQEgsY+53
y0Maid9HxBbWMhCmQ5TOVN/tCOySnshwOGj4fknHaUc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1920)
0o3B5IUyPNHZHjWD14iPtNrsk+ZN9EYggnr3qt9fwaF/9wkSHmjNGG9b0WfTQg8T
WSUCDOHhVByyaWSw6RyOdQ9uHodg9P0oU/VAOtAZ9S1mISZHPtXtnjaTCGCmrxEQ
slmu71kvw5m+rPFlX2if0ezdSK8XipZ2HBz9K4xB/5vGqE+R2qe588b4lmo7a65o
dvMMXPPo2gqVr5pGdJsQ6EsNZaW0iL2yhcmt9RIBB5MXl+GtKa0z2h9uAO7HIYUi
6+OfuTIaOLpJhrHyyb2r42WsqRmLdSFbTz5N1gIHFbq13g2bIBYBWcW+ze/XirOG
COQGLda8veUqRC31EayMIck5YSMN/WEq46mIyYm9MYUjQG2NPpiFAg/Cdrj/ZRdp
hrXMM85FIUdMrjGSqkG/hq+X3jUZllQWmOJVULyehTAaqL/Ogm8j0xQHeY0P7/5t
TDWa8Kxs9806LpVZE2fDkNIGJ1oQfqpgsrOa/mgGY2E6GxrvMNw+X8pRMCIYtr7h
aLJUy8apcipNyr58eebQPN0jG0RsVb+QysHCGJngXWmnj5m6ovu0+RBNnDS6+nsa
DyDhu9mqe9qyVGi4zt0AIpHImOPv+1DwO5Bk/L5aYLGggKBoiJJzeVTi+Q+5ila7
bwfY5RWhdXm2tSY2mtekyLAGYbQZMTwzYf6rsw3Hxu7zEb/WhyLNe5JWCBHuwmB8
8ljDU4vEwzzi3scXZdvuDR+c98/Q/5BW8KwBlhJGG5NihdJwybmjSHkMt525EB/k
sW1WNrgfd3hM4Yuxvzm0acOyUPvUcu5Hn4RzGiIRee0VXMIQQ2CZCp/j3+tKYv0/
C1GkYxqIRMFSl94956RGn9IadPWWY2N7HWR6E+P4XwAGSCG73VFkYkIBWxxXQvEJ
hz3lrt27BEfRfYugAMP43aT0GjVX1C+1TmK/15A79MteEqRNcBm8fOmxtJPTcN9w
4xuHSVIsR9D5IORi8a3bIxEGk9e3/g5Z1ByPFvSUoWVYiGwUnxxq+l6micledeiL
h6z6Pormus47AqluESeu/+L+qTuNDoIkSvPf/gkDbkHtxS0kiDPJ6h8nmzzqejzk
naHhyurNy2DJMQ8Bxm4QZTfpW3HBlpynA6+bFUQLi6y76YKrR+4c4MVhlxxNweAP
T9zxV4J4zV0Zr6Q7VWOEJZQfYXRTEpK2KcIO37DXz8YIKE+PrQid5BxYhVVA6f0T
fIvd+CcniW6p8xftkv7B/u6Fo9JNpDFDmiLX4cxqaYw5ZHwakTICrbEH8pPODH21
xNE+/XzUtiTxQhsvQkxQ+i4ASdcFbLmaSql4wuixabvQjWjHtSGhVCKMePWR68G2
38mTtDY0HT+xlXG9BJA95zTUcOiE/1WuCJWbvMvUrMZ0jygJMvQbGR3APVwcR8Vl
Th7DDd3oR/kvZCIkLX92X4kCQV3bUCh3BfBpUnroj4rIoBwuNsQSpgc76YQH54sk
1yguHD+Frw0/JVI/xVqCpT7jIWk+P913DVR65L8ZTK97y0UHM8Ho236H3jPZlqIg
fW3hQVSCYc+03HGaiOV+7II2zklx2Hg/XTXMkGGbql3ORkLbjnyUGhTOEIpBKSoD
6la1N1qXW3+syRXn5q+W80lKrUHZHsiyrEuY9StTRIAU9m5Hum+ccrSHJaxD193y
nQrskSls6zF1WBlNrrNYcfG+u941/9wqYvSJ3EOQNsTb7mHG6PQQ+l8JkiExvdbz
pJuNN+LKIOQ8mqvFZirK/kE3syCmVvp03+MVai0qOQsSkkZeNOHtfLB7NoZMj4K7
YfanDufNxk3QfNYjBs9u0RU6JS21h1VFUj1jFKKHPaj55Vm0Ua5rxnIC1bhWi7F7
d9NuKnK60vtsYX/90YQki3HYh1AnXZofLGnrgUHrN9z4ErWyzzFr/OFg+AYvwC3B
shVqMmcqN9M7WEV53JLIncrdbHPH+QKdZUwOrEe0kfwsxZQzIBQu+t9goc65bwi8
a660bG/GwajAAZzyjtS0XqF9WEz8WTRBvHiMI3CqJzkzhOTU8BEarRBpvHHjTDTr
KW6DHC0GGWZHCf5qCTvJkU0HmXswjSAt7GADbH8UqfA8Hp4ddgWy4aLKN9eDWEZ+
1+Ia6Kax8yss0OAv5aqhs8DnzRZzcjfSXCIQ94Y7W6lsJ2q4kJZmZUcjG2zzrtRU
GawGVYvpcSOpkIvscDSowvWbe3p0BJOM3mSrJs4qfTkbxVP1ZlRYy8NsXpYpehGH
rxkFr7eS4Ooo9AAzpWqEJyFH8SlsyS+ihZ773KIKc7EhDPp+PMQYNHL2OzLbdzKV
/Wrj1Md3u00y2vsrSa1NEGQq7dGt/M+huEc4j/lP5cqaKSiClSaDPDDSivqckbi5
7hkiDL1t5STrVyJxP7UTq4QaHdheeJmnfftpyM7pW7IjSKJfX3PlEExZMp9eORgG
082vM7Q7UBz9GIpt3Qh0YgGbG8zpxaXUVayP1sEkJyuUjxU7TUdambuc3Y4u6OnO
Q7+KIx8vgC1FoPsYnY8SQKXGQPNtM/cq3hv5U0N0jFLjMrlC2NZCmqMEmLSQvrCl
`pragma protect end_protected
