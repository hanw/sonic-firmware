��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z��ҫ��=��� p!x��&[K��1��Td� ��������!��/ןz��z�i�۹#��9J�/uN��g|�D�]@I�t��@�� �z+x���R-(������@����,|6Y�6k�'�X�W����u��=�}��r]��n�%ˏ/�gr���)�����:� ;"���;�}�O($���M����;dFt̺�Sey���P����f�k<��{���/�#����?�~�6�r��خ�B���͜8&�;�� ǰ��̈J�k_`��]�`�拃�R5��P�]��
��N����Y,g�UŌ��`O��}y�����Y��^��B���!�7��7т�U��"�B���5ql6�W�8������2�|G�(>?=O�
�(���_.
��S%�6�
$!Xp��(ŝy>�D΀k�1_Ks��(ŵ��p��7����$��
�F�*��%��o��*1�Jsߑ�}񗬤o`ZC��L��	j��Z.�� �e�&(�k6`�v͓~�J���ce}`F�`��r̖Q3P.R�阮I�H�MX��j�)��[�(���'2ԯ�`ipg���������#�A�5�1�}%�0�u���C��#�Yׇ=�r�2�W�.6I�W�c��pR�?�g�Er�ą"l��Pބ������������O�l��5�|o���;0�-�9��$D4N�M��+���/^}�*���&���%a�zE~���a��24�Vn�;<-k�w}	�}�-�Pi6�:׌���_Y)T�Q�dm6��M��q���u�Қ7C�'/���*��0�Q�[��wc�Z��74F�	�U1�e�H&ݍVO����/s�BC���$�J�y�K�P!������G)��ɳ/�"��e�p���[�[Yh��nGEDp��o�����^Z���C���H;_v�r*"�(�44C{X�xx�ٲ�����6��kAs{
�������\�����'�~�<r���Lmz^��	A�/-��VG��#�O���h{�͟)�i�kS��
P}��̊<�]C��	y�7�6e��F�Y���A��*]��l��x��9D�tbu�u7?�O0���.f/XI��D8b�v�}�����ɗ�r]i^Q�)D"o�_�2�S>��W`��ә{R�oGy�Rk{�t�cD������_�MT�C��:pۊZ�x7^	��ʝ[�����fE�b���%�#����S��pa�-C��`��Ǻ�"en	��\e5M_�p�Z;�O���@`� �οI6�$����|�EN�k�7�3�Jk!i����ZԆ#��}���A�ׄwQx�~9U�f_	���R���bk�+�o���E@��d���`�pR���i��5Ʈ�b����?ߥP֝��>��T�J�x���bѐ�!���>̎0;��Ļ�|bm�V�!��V�sC���H�|!��S����\?��R��m)�f�F{�;I=C�cv����r�0�%5�%c#Ha�0q�T*Չ@/m�U���A���Z�~��_m��L=����4��XR����=����@s�aG���,j9�_Ԁi�쪘Y�XO�;����g�'%�\[a"qZ��9��h%׼���;�i��!��'A�˔�D���ӄ+�YdH?�،F`y�:]cH5�������a4�b�'�@�z��1�9��N��i%.CҢ�I�4�XT~Db�;���vp�c��,�(�z$�����i�Uʓ�,�f]����|���鿍��E+�U���x��D�:�I�\�2�ع)xG�vf_��Nn��%��Obw<N��j���n̼�|��`��N\�<(��*���%䖔M�^�B8S�(X����w�4��~?,G 7!���Q��/#VRyXi n��������@���[k���H�:��0MZW�3���DˌE>^f�$6�����ܘ�H��9ю.(z�!lٶhC�h?����N�"1�]�J,m�"^�A��_��YZ�|D9���:fp2v1�b��L��`�((X���<�)��P3�'=�*���ͪ9G�TY����j<��G�Y�QG��Փ=�*s!V��i_��qb c��Ç���ӵ�5j(u���W#�扣*?��c1(]t�_+v�.��Yc����5Dʝ��������8������1Ã�'c�m�R�PUE��V��D��~fD���*:���������5DG@V�B����mYHK��&;G�Hb���s�?�u7-�e$9����e� �-���{���B���2���p#z�ϭW� ���2�YԩiwiM�d5W�y�5 C�@��g@*(p6j���0[�|x��xTe;����.ac���e=��E.Rʤ}����0��;�p�X�������y�me��&Ut��n�kː�)�K�TT7x`y��r�,�y�ƺQ��K��7�O�-�-��ƪwM��3�0|w`��l�q�2�/߆��d��IA��͈�МbܗpOXN�B,%(I����ߒɛ��<�nVΛ���h������!섟�3]���꾙������0&�z����7��L��X����=�o�-�:A����;"Jɹ���
,xf��H�3�%�������(LB�x�۪U7�s{_Y�[_z̔��C�ͮ����!�7��u��*�G>-G��UmF��Fr���hU�9+Ox�-e����~�5�SVGs���W�;�:��d�ނ5v��$�2�|i��o7��?5C����4VV���Lѯa��S @TK[h`М���SϺ�
�~�oöq0mX��y��Kc�ŬwV���O>���k�`8�3�^WK ف�P�S��/��M�^/LX��U��Yi�/�����,�^�����0d�V�M�\#[��_t�Qo�qH=�х���6���L��[��Â��h���o`(�����Y���0t�F�4XMA�#�)T�M��j�8���f���=I4����@V�n9g��� �8�9J�cɖR��̉U��}�BP�:A,�ZeG�����	���4���2��ZF���;����#
�NEv�t�w��)�;ov9��p#�T����Y����XK�bi����]h�C]�� �T��E�:#,��*�����-U�Q�� s{����~�C���A��,P{���[����Y�@g��%�|&KN��]\����۳�y9F��ԓ�%�dlP�=��`?�K���M�5�����i<?$i
f�y� ��?)��e��]&�0�*;Q?�|\Y�x�����i��'�νR���"1`@!F�{n��G=f�[I�,��UH��7����r����ƻtw��]Rs���|3{�W�FO�Yn4�\�ʭkaЌGL�1ٛ%��Ψl�Lq7O1ԍ�D�$��+�����I2�!!�h�g_;�|�ֹ楌6�'���M�F�ll���`{܆;ȥei�SwU�HҢ��c4"+
��.�M)���<����tUO"L���<��� �� z��n���P�>�U��n�o����e�g�ms���Ni+`m\N>a�@��s\���;3}k�g��̲�1��E�*�i�~��7�>�s�wxX�ʱ1b��捉b:��KՎkF5��5���\�\9|-�Np�#b�m���BjN��\���o��Wb0~�b����[	���Q/�6�v&�$���������+a�.�wn���'SgM�t�ەbk�V3�ZJ��M,#�k�K0���L�/�+�5����ց�o�A�z"#y��"~mN@0	����
Zת��H�Ȥ��b�n�;�G�c�"7��}IX��cr�j����p�L�贱taaq�T�#
,[	��Q���7^�c�b���J��[92��-��-��:$�S���xv[1
�<N�~'W�s�Lc�ڴl㸗ja_)/Ϧ皫`����0�P<U�"��D���<I7����2o��-�֢�:�9�)��F������h�������a6f*�c
u�W?��c}��t�M�溜	��VϿ���V��2v�țG�Z��JI��9N��u�F5<y��R!��3/�/�Pj�}����V����
�{ml"M��N��`o1�$m�lN�6
�_�?��$%5�5W�,ZK�f�Vz���>8$�_�;CQ4���%c�\t�$˖:��"}�g�J6��l��^/�>�ˢC���v!D�h���������F3�`t���O�諾l<�Vq7D�#�D��B�e~��jD��M]�?�!kP�A�|�RP�LSv ���}'��#�B�݈����@�|��ΐL�������'Z��%��5���.#�4m����N���O؋=,�&�ʮ�1|�"@1�nO_.7��d��w�r��OP�t�G�~���iQ�����(s�ry��3-iDHH������3���:���U��b1"�βl&�?�t�,��Ha}��+�E0��R��%�vg�����a��cd��6�tiI��JM�r�����dC���]�C�PP��(r���G���|�X���)�߹l�
&Th�
�Ҍ�kj��r�\	@����^fS/>�xr��Rd���o�߷u���j*$N4�Ip�j���bl�P�V�߸�>����5Ne7��h��>�0��9��#�+ks�pwݩ���|A^�Z6��7݄%�CG�$�
(�ݠ�[\��/��JY{�FnU��Ql���d�E���1�s�@��q�Æ⵲�9M��Vt������|#� ��H�u��¯��Dj}Bo݌��v��f��c�sdq����W��%L$ހ��]J����Ql�)��9	�$T0�Z��K!+�6[Pi�tY��D*��!�U1Mk@�[``.C����`~L�g ���9�S����u~�哂��t�y��j�u&��o�^��ѽ貞�T`�O� ��Q��v�G���L�x|�Y�Zb�D˜��{��"]w�in>�΀��I^h�������UY�pk���&r�|F��xl���C����A��<�I��6Rr�d��n+O��:UԚ�F��tŅ�Ctg��u��-{0o��Jf�h�>yA���0�@�D㥉<�+"ٔ��Wx�H*c^^:�����\OP2��aP�^��}�i����u:ʹ7�"�S+t�(A��	�i޻x�qNܐ��x�Yo�5u2��,�CI{�*sxK�
~u:�����Ѯx��Z��@.z5�oa�؀����C�y,P���v�Id��$/�zg��#�����kwg�1+e-�QrmC���x����䋨z����kY��w��fPd��	��(aɵ����8��p6/���7ś �L��L�H�v%C�̓\�.�\��z,.��~��]�7Q��y�J��j'}�yC���t�B�0_[�bYT��9f�YN�ue�<D�����S�@��܈HT�c��*ͥhܑ�����}��I �ֽ�ʖU^���in��p��.�L�<'�����ĒݦL�Y�}X-��'_E����Ǌ.:�rjv'����ᗘ�R���Mr�4����*�R?������G]·H��3��w?�w��z�Ȼf����#v2U_���� � ��-���t�����?^���S�K�����	.������VRiSk��Ά��t�3m�_���V)6��j'�aH�����^�B0AM%�낋qH'�O��嬁�V[��.%C��5���7���Ir�ɩt�M��A��N��� ��S�Om��F �.��|�հ���l�G�y��r�+Ko��V鶫n��׳�v�U�ð������'�3U��2�f�pT9Č�/��R��9�����׌h�]�h�������	�֧�MDYGs�,y����
��U��UgԒ�9��:��x����t!H�	^ l���
G�a�7׻��g:#��!W�:d��.p���S�"c�I[�K�'��7�͗>i�����b?G���H�}��E28���UQ�>$-�P�H�hs�g�(o+�;��������$|��,�VR@Q�K30�(�#eա����Y���	et�Z�>I��66�=�m4%�s����[�)0Vo��hl����:�WS��>,�\�H�q�ί�H~��>�*��<�����������^�إ��1Ykj�hD~�<�N�6��޴�x�L�>�=$���?W�S������i6�/P �0��.A�k�ByC FS����W�6�c5L�R�A�u˺"�aǓW���H)��qǉ
�E���+�c`�7�����\M��./�;��u��:�m�~&q��RY����lSȺ۠CX�$���At(�5�qk��f6���(�C0�m�y����\�K`������W���ɱ��f�#'�W�0�<��$�}y�0�� x�W���>N�h	�_�ܬㆪ	��u�. �Z�N]A���A���k=9�z��ߖ�ҁ2���+���p3�v�8���Dz6w�s8��o����Vy��	��ObB��ԻEWg�K/�`�%d(V���{�q�y�a�ԫgr�%@��4q����$��u��qWH�BQ��Ҭ袎�h�B�X�m����Q�[B�D����{��N��g T8Y�g��p�����t���	�kGg�܉zOS{��<�39�L�Ծ6� �8侪�x�d���wֿH~.�� �,O�@m70�?8�^����b�ی�t���N6�Q�����>d.%�'hs��*��/�P$t�s����_2�hV�Z�~��~r_�KS	ը�1ʼ�f�!h�W���U�����Zʖh�/�ʻhG�E~����)B+��CJ��W̱�e�4wR+�-���R��8�����G2F���b>,m�u�}ϻ���A��0h(~:9bD2R����><�I��#j� ��G���@q�����8P^%na�&�^\�i�bFK�22��Y{���yQ��Rpf���7&"cj��Ei�&�˄�f0�r4�qv�R��i;obE������bA�䕘'�ù�ik��P�j1��9R�;2&&����IS�r�����K9���F�Hx�|�L��w�v���%�,"�5[F������F��ճ^�m�i���^G�Hj��myt���������?�����w8�_�9j�8�{Z�::�v�*������l��#/N�9f���#:#ŝ�/����WvݐSe~V	��H�6݆O�`�Æ�ĽU�9Q&ݹn$-�f�rU0��3>��R�S��Yd�k9O�?95w���2lW�=����澋5�\�B��C�KSb��ދ�[�i�G�q͵|�h�g��[��UX���t!�l0ݼ��h�g�ܖw�,ݫ:�P�~�_D��������ʬ�Qn � &�&���6 s.�u������?���������N��ѽ�Cgnݠc`%�9�� v��T��sH��޳���������
�?7UԴ�3��pe�@9�8vYK-��Օ9!F�*��(�O��oܔ_�Yn	}���O��"�:0��Jcs?9}�����ڔΑ#wN!�ް4�=4�[P�CW��JW ���&+!�t����f�Tnka[�����.%�.<G�U+)8<`[53�<o*����<+;?��/�G��.#2�^,���9�=E��>G��s�!���嶩P�n�l�Rp�>Z�{�ƱE�y�1�&7��3O�D������} ����<���������t�k�hA5��ߥ)<�7u����4J\m'_cxOk��U;�
�H�A����Q��Q�����T�hw��^�K��
-d�p¬�ĩ+�����'���fZ�j����4��G޹M�R�{Yp��҅$K����d~��7�ٝWJ���f� ��S*��p��k���O������o1������)��.|$��&De�ŋ��*�,xC3��L�(�H P��t�fl�њ�I%�>*ԋ��=�ث,LV�1~���T{@���/�,���*��p+��/$D�N����6"֚Qy����/��5��@�sno�M~,��Wru�|��:" {��uM+O��l�����K��"4�yg��@���������ʪ��6r��l$��Cfbx�"�T�\�d�%@	؎GN	bd(|'!b���[AP9��^�q��z������� )|�+lJ�nqO�N����x2�ɧ�`N��j,m����ݍDyb�#�|��i�������� 6��ɏ��A{���^�8���[}�<eEf2�r3�,�S�x�6��qʨ����g4���0��\S{#(	�eض��cy�-��,V�5s ���6���g��:����Pĉ#�Az��lG)��_�7�r%<$�Ƅ���Q��}��;��O�cG����o�=b��J�H�>5��ԻR�Kv$
�v 9�K�/#�V�}�,J
֊��v/��ϫr�@�����c$l�,��#� #,#ՍiYJ�˥ڎw�k�Y��J�r��X4?@s�0q��Z\Ĥ���uSa*Vu���R���]f�?���wQ ���H��	C�8�#���Nbw��.�O��ѽn�uWA��9�Q�y�3JD&G6�W)h�^�V�{���)�w?i})]��
+����]Q.���f��H�嫅�"���%ThNWߙWi��*�ӛ���T
���cF����rk�̫�y�L�Q�GW�5�uM�:�����]��K�Ba�M.X�~�N�i�i.��fZv ���h��H�l?��.���__Iv 薮�W@��w�xJ#�qo��]�a|5�%�+��k�k�Z.��F������2��8%[AKB��,���g:��{蔲�Fp��9�L�q��H�E����t.�w#<MeB��o��z����g������!��V�{�Ѱ�viލt��U����7R�\f�Y#�y�oR#��F�*':��MU�C���Pﷃ*վ�<q�Κ����
��8���Z�V Z�M�zRo&���ۡ��;���?�� ��^��Ej��A��yMh��I:�.�69�#qT�S���B@E0�hoN��9l�r�q�ϭ�����=�Wp�wy��ȵ�b�w�����^m �����`��b�Pf��ؾؿj=�.f�<OY�f�O�4��@ U��T�U��'VR�b���8�{�o���0>��"U��n��)��z��n���?���@\��g�}��K�ݑ��b�r����(�mͿ��Oy�j�C�ѳ���L׽��fP���
SuR���5��c�$mnu�>�VHD!�|��m}��e#����֫�W���	V杛��{N���TM
R�����k&�|���d��ֺޣ\���p��Z��XF�}$cf8��H���)�bU���tcb�mZ�j�v�Z��\8Wy����٣�&k���}�h�n ��W�uf�y2l@����a|}�1��x�B�:���Oe!ݵ��=G,?Ut߽]�T�q��腷F"��a8�A�^�J�X�	D��$#�9�KAⶲ���U@�������|NTr�+��'Xa�WP,� !���Gq�r� I���v���h=G�����-���b�ؑy]�{М��
;��MmakU�m$�����&�R�Xb�EB��	@1-�L�i���Ey�x��{5!��BbI�E����(ۥh��^��-�g���.�!l)C�M�Q1�z�J��;�ԙ6���@ T���6���N�9?d��/��C]L(�Cf�9�+���k��ʻdI<��+%��"ȁ�iF�AO��V\���RˏqM�9T톴+�4��H3�;�,\�^b$�@2gi���ډJ��>����8^fb�\|$�j�VKgN�x??������`T����%al�E���=0Gl�������0���[A�uq�����, J��EϐzR�Ȯ-?�,��׉k�PJ��9��G����䯷KP��j��bOÉ� a&6>+�lj�f������;��H;�q�9f��9��6r�%d��B���i��ݸ���ڪ�������t>BX����jKA�O↲4xA�5	�l"��싫4����A_d�j_��E�V�Eor��F�g=�p����9��nڃ�����3[N��l�эL�;x�x2�������&�R�p�MǊ����7�d�Nj�B�>˩!�N�������!$Π�ӻ��8����(�j:�������D���a߬pa����o)������#'4!y4SQQ����f𐏧"On���8���
q��_�p���`A��kd���w7A�Q��J/K*,�8����&�{���a  �&Zx�I���[Ƶ]�Kꄂ�G���5 �P(G߸5�紓lj� =r7@6#���B���tE;�G@1���E@.�5ZH�e�~s���7Z���!,o�}q�=B_�Ù�x��a����e�@	�T<����d��>�M�7=��	�	���4���@OA�R��4�о:k���W8Y���!���%�'`�9` �1 KO��(p��?
|��N��'����׌z���h �.;Cz׍Zϕ�xz��=V��u�x'�Մ�rOjZ��/�TW�;ٸ��$��F*�W���Ϧ�>o.�A�k3N<��y��,͎u�М�&�֛w#�Q���'|E6��Dm�S�Tp\�~<.�wX���L�2A���Mt%DД����_H�d���剡�Œ$CC�>�4�P-=��r��g�ad�g����|% �o���j�w|����(�vh8�mA�gf�0c����]�+7�y���wī��H́)t(��T�~4�A:���[���OA�>E�qeh�� �:��<4���´Rɫ�D!�{���f2�`���#x�"h+B�P�L���ezy��޺�W�b�ܹ�r�6��A�䪫��>tB��"d�m�-�
��o|��P�w��h��4���������i?�Ӫ��gi7RrLwF�pT�o�P'����=r[[�X5�� m�ñ�����E��U�6� J�0�trs n[Ά�����C9}��٫�h�M���T�Z�[�nW&�>��n��5ϯS�3I*����%s���������>PD>mch�0�]f���(E��;�F��@����N�+nX7F�k��X�.���T��L���|,�����s!��-���jW�n�a��@u:��� ��q [���U�'��碵��ͮ��J1sZ�~�s�j��ܫ�P�N[Ċ�N�8YݸIb��rɚ~��J��|H
�����ب���@�&��B�~�_(R��g����z(�nu���u̡)�f��*�5���$�Q3\������e?A*A�8�LH��7��ٚs��d���鱄h���b��<��] R�i���w"���_��{j���]�wk#�%���[�\�����d4��Z���a+vM�kq�`��.��fj��{n�*�]�������\�Zr�e�&�����|��o6BFAGYFeS��٢px�E���x"�^�B�iD���W�cE�Qt*��ܜ��+6�ɏS�R���ut�9.߲��h����
UCC��4D}�T�7����	I��	 �'ޞ�2E3��{����1�[��WH��Bq���.Eո�tIo�0�Nm��Z��
TuNg?#��'�aG��H��f�u���T�V�����5�4�,Y�Sj�1�}j4�N˾�I"�RU$��
�-�exzrDwZJ'�<͈%�h�q� )�:�,Cl�AQ�F�2v�
|������Z�
~�kXc�CdYO�ɾk���/��4V���PW2�rA�=F�s��1�R@�WN����~o�Q�8���|}�қ��	yk���5L&���V���sG�TPm�o�,��y��sp�m{4�$?��Ɔ�~L���J*�ͼׅm�R?UG]���4�вPo���wI(�;�m�K�$����*�$�'��+��O�W^a�D(	��Ϭ��|x$���|LI�vݗ�ec�6���v��2�c�����a�V}]Ѫ^�
@����ы�o��$��9�s �S�&�9�s3:�����Y���M�r�1�yۘa4E��n�X���w}�{���^��D�\e���Vj���v�����h̸�O5�m"�?��;���,���B
��`<|���[�W���x<26�2;�*h*z;�q��6z8��Pr!�E��N�^w���ä�5� G��w����_C���7��Ӌ�!��7����_c��Q� ��H� 9�-u��8���$�'�\
@�����:1[X����SQ��ΞN:�_�e[����y���giTӿ�a4c�r|O8�5��ګ�&0���3���׿"�Pv�c(ҝU�����W(���cI����Эl��Q��i�m���/��ʵ(Uؚ+��.�P[��(�d�j��k��4�O7�49� l�~��)�L?W߰]��M���i��z�qNwפc웉�--;�?�x�Go�S~%��
T�&�7�N#5�P+�:�53�B��6�˞�H�o����"|:XN804�1#����ӰE6c
~���*�|yABm;Mk-����X �X��R��o�����o�t쩥�s��N2�$���톶]2�7��]�_��i+x��]��9�:�.Yym���ͅ����ז)ʦ���&�y�L+_��������83۫�<G)��]o[rݣ��z�_�*�=�/!���K뿸�2K�&���Y�� 6���>I?^��OQ#�֨�:-��G4���8%�cf_��〔���8Y�*��ϡ� "O�B���[��DR��n��!o a�����ƿ���)5a�JnjC���p�W@Ӄ�D�QM3ivL��0f�"��^rġ�EDa��b�	�`�u�(�¤���m�po~(�}4�������2���q}�EU�"$K�h$��#�7�EN-�e��ro�nXD��D^����==IByqG�T a%�`�f���5o���<��.G�A]�D�������h��e�!��'#^�F����9�q�wb��F~���Z��-T!�x$��3���r���٢2z�K��<����mm��f|ŖgMڋ�γ-�#V�)l�r���������TibL R�a�5�"L�ؾ�9l<��(��!�=�
�e��j������х$�k�B��A�<�<#���7T/���'D��J��.�B�j�v78>��ԯ��B�����f2��y�Gyr�v�����V-�<��5i#�u1�:p��OF=�.8�
K#.����x�޾7�Kz?���KG�upI�I<L*�pf{uT���R��DV�]񒽍X�!ʯCx2ŉ�5�7���uL�&��T+qW= n�f���g1K�9#b݊!GB(��~57�X����Gc�_/ܬ��{�����8�&�!\*3X.eW;�!4#��WWP_�O�cq9�[��ź[=��v��+��J�,�z��`���:Uo�w�S��
;���V�jV� a�[�3؆�V�c��2��	q�6H�F!6��2��_��g'ˏj%�~�=K�Z�h�@������ss�o�s8��d��kbd�%mS���vOכj��8s��wf��F��FՖ��Ȕ.�(�����3�b&�ZOҾ��ݕZ,!����p��0�&��������\�iY�|0v�ݍ`�K@��i���9���'�������Ofs��w�=���Z�y��r��C#�hQXΚpJ��Ɗd=�1�ۚO�1�g-sL� KkGz�bOg� �O�]q21�jg^nZ!˧!u�I')�l�p|<�I9ɗU�;�V���wB���x����u#	��&w��NY�?��媢]Ƥ|���K9���;�o#FuSf�/��{Ga5���䣾� "َk�+�3*����'�]�m
\�GJ�37Qg!�-������L'���>N�9_|�W©�Zf:)7,c�p�[\���Y�}�� Ӯ6���C�����̭E*˷�L��K��ĸ=g��5����!T���Bv*��n�=�G�.���hr?2E50F���QG��^�����-�4���%�懆_zi��tZ����� ږ����5Xׁ�?Ą#2��c��m�ڎ?�����q}qތm#1�0%�[a�uo���zۯ\��(>����-֑�7��8l�����IP��0��<�:��������S�I�K�ӣ���l��9%(��i�l�\ppt�,� j�UԚ����r4e��*w�E�h0x��S�����*���6�`���I��n�ͯ��_
��8�CZkz�Eɚ�*�?�m��hOT}wR���U�����_Ў1��p�����Z� ���n��Ӫ=������m��*%H�{#6�'�����x�S�`��������J'9���vS��O��8om�"�`��6I�Nɥ��g�V&g�΄|%H�X*�sS�&�O�oQ2��tpR��r8��Z�1SD�+!u�o�-���9��I8��o���)��
eբz���ԫ��5��D�=�l��Lo�hL��d�ݷ�ᐞe�Z����t)��A���n͌6�0�.��dRz�3jk��.�0qГm�RQ�H,�ed%
A��$�����
*�<!m�2G�����#��x���ڌ.�p�w�K`u]KRka�Ĉ
ϊ�D�"���A���UpŖ^�?2< �J�'($MA��=+
i�|�p����?D�����dZL�(!��R� ���]�L��48`۽RmS2�,$v@5��,LC���n"�����5�Sm��Y��f63�॑��[��������q�>�蒠��f�J@�8�5@R~��Out Nf��p�?���|��K�r�on���qYr�l�.���ƻǨ<����!2�P��?r�,_��jV������hb��-�e��M#�Ig5`T�́��/�-��$I)���ʹ�Sb_�'N�,�H�S�rƴ1	u��z5�T�$f}lb��z�5qg���ɮ�w9��ZU�|�a�zlǙp�C�0�L�!`��@῞+]HT!�Z���f+��j�AEqצꌑk��r��j�fy
�H�U�lK��w�,R\��bl(�mm/�^1U����g|�ep��͹q���m�ZI��S���K���c{���Ю{f�� %
XI(�M~�G.�K&�M�'����PC?�J%@��6�1��x��C�s�8�1&��q��U]�	�_��� �	�ˎ�w���o7������.xtg9!��Wo~�^��1ؼ�.H/-�6���mG�	eF�	��Ka�%^P.f�YX�&@!��y�|�=l�'�Xa�����>�`�$���^P1=C�R��-J�<�f���*���ٺ��j�Y8쑵_t����Y�z��w���*���d#���X�p���KO���t��z�����Y�L�6>۩�|0?O�O�y�]�9�������j{��D�:��t�5�֯�IV`3!|�W 6i{}+b�W{ȜNx����d�H�������vHw+�H��o�B�jӝ���Bi�-��Z�Ӏ�YS�����8kr��e���v��|]�9�&�:X�3�~���Cv��D���#�2�׸�