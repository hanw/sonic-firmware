��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z���+4eTc��� /�TU='t��~��S�=��<��{5� ��4�H�t<��L����z�`���=��X�L���";q�Ϣ`bk�aڹy|��M�0�>���Va�ɫ������0�����)���d��̸Mn��-�r�N
�|~o�P�Jql�Yr��<��"�:e+��/��4F�X*��k��G��Z��V:���`b�g�QxK|{�q ���oȺ�BFR�����m�9Bv��6��1��r�Z~{ �S���ݛ�U��,B��
c܀'ɀ@�u�o򐨕/��Ԭ>�7:)3�vyg��t�מ��g�0��������$wKd��%	��o�Pm�oj˅��fl�Ȟ�a�}�n�Xvq!ث#�,IB���z˛*�r6#Žؓ�[%w-��g��H�hܩrE6�}�h��zF��[G�3ˮ#.{�w!�Y�TǛ��m�B��쑒�0��Z�[e+(�1!M���h��i���d+8��1O��t5s�B-Ͽ��CP/�����"숛�����.㏣V5�j0�DD�շB?3=��l�l���<n��c�������|�ӎL����X{��j	���.��s7���ґ΅�Iϔ�E]�r��_�����c�c��Un��ml��ZR!�C�ר���`�Ź��Y�^vM�H{����tȈ�`���_�;gS�p1=�/��F�|"�F�p>��_r�%��?�e����2��f�P�͔��q
�f�kf�I U̂.�L˸����g;�وn���H�x�O��l�E���5����U�,�c�ĉ���7 %s v,�Fxbf�_���W��l(��_���&�v	�*QTЏ7q͚�%��%s0X($`~P�ˈ�r	}�����+ۼ���U�p��^�D5�E���(�I���M馲 {���0���~r_�ރ&����=3��z�������7�!��]�+Z�3�n� �r4���z.��^uf]7���K�2^��F��(�Jⷓ�c�u^M�0�@�/�hה�|���=
�0�m<��XX�Plٞj'>�vb���ec_��c�c��ن�x�s�JS
r~���^oD?x�T<��\�q��%]�Ͷ^��K`��u�\lmf����ou�K���wwX.{��61���&>��
���U�Y X�X�7ZX���s\��d�9PЧ�u<I�Cҍ�6�)��Ռ�		Յ������s�yߒ5r.c����]e�:���R6�N�0���v�s+�]�>}q��Z�Cg�羯��G� �]���d�]��Xpv-pf������'�k)����J���b��f�9/иNz�/ڷu32gt��Dl��Ö�M�yJ�c�T�?��n��>N� �_����6��s�6���.���<V�V*���SٽX�uZ{R�b�[N��v�I�_VF�
��ܲ���v���y\~e�V\��@�u��
-,��D-Y�^��>�u�?W�����<��=�)؟$7+^�f���>UF,��3�)r�h"�.L6 �ܱ�ܓ�{�R։�G��#�s�Ж&T��X��J�Ѧ؋kQ�a�IN]�E7eԳ��F�$q�V;P8|=j0?zg]F�{o\�8a��e*��_�tP<���:����ssN������7���׵�󥀺(����pR��L!����g�O��������3T��X��s��?��5+I���"��M���̽�q��U}d������A�OD��҄bg݊~�%���:�,�,N�e)@��ꄞ_��,=►�-��86�(���Q��~O��r)9�P��C��X��ѻc��N�-��C��γ$�f	ʰ=�H�JSt�c�����L�_�f�H��H��H~��VT�����%��fnؾC�*bN%T*��` c�\��d�<�^Lխ�atp�ݮZ�.�J�!��׷q�C����@�A�)��W��.��oW��e���ԫ����$���]�5�n�,�j4�kh��!�K�"�_0�U��� �x��̉3oB`M=mM��� <�x�Tm�0�[�R�޼�Hc'=|6f%�o�-
�G�n�c!�c��g
W_���&r���3��-���hQ�� �m=�f;D�9��wF�šd�ȵ�휡)?鹞�7W��b�u�ĭCV� ��2�CN�X�pڔu��v�|��ʳ�Fa/�17���0T�[D�[�FZ�8���7��,�+*�_��k��fӭ���2���Xl�����3�-u�FJ��MkK]���C�l��/�2Zm�t�MO��5@���L��g(^e&���-%��o;�%�PA.X^;��b����)J�ʴ���K��@��0��{����{L�J�9���k���$ټ�.���2����FL�K`\%jW�:^L=�O��JU�]#4⑊�u%��7��,�����Tt�'�����M�d�׽��8`8e>Z"��Lb���6�����?Hq�Ɔ"�a�����@,���L�mM�Y�� �N-b�8��'�f��Kک�լ^aU�J;�+�c$�=)�'�Юr��zM&��F��K��c��A領��T�����m����u')� \>���
���Z!�B7��bft9Ws�|ӕ	&��%$�� !o��eM����!���쿸|�|ޕ�`�y�������C�	�i ���s9��Fe��M�^x�A�&��y�C���
nA�6�����]��ve�$Y��O�f�<�H幧���LW��ĕk�P�Ærwj�+��c��	7d�P�ܗY(��Kj*
a9&=�HL�긕���Zb a2����0���V2k.+=w|j8�"��B��p���6p��w�6�|!g�e~���`��;�^0��)�"V�U#��ۍc̓+����e�Fc�!���G���4�G���?N�-�ᣬ=����8�����w�]�c��`ZH9e�Q��2�} �7
�L���_��w�0�5A�x��n���㭙4�F�b%ꈲ(e�+���؏�'͹�*�K%�=w�L\,�������ݠ�أ���LC˱C�->֌p��X�L7��g�E"����O��ݒ�z�� ����2�� �ٱf�5��m��2�7V6�:ګ_�ܪ�6� ����ٴGRI��_!�h3^�A�����'����3���c�q5��ӈ��O�����%�i.VP���=��or�ϛ)ȜD�`�L�
��8� ���;�~�f��p.&*���a;\#!)DO�+]%��{Z# VnU�W�:O������v����R�p*t��ɒl���i�a�χ� �� �U[5�<lvE�5d_�J�*Ċ��=VjA��Y���oa�6���:�}]<� ��4q8�P�p^��\��,/�[	'��^�D��6�w�����J��8�%��q;-y*}�2�l1�m��N�-,����ä�C<	���D8��ʱÓ� �)��z�lk]�j ��=s!�ڲ��*o"�ae57�<yI�����=U%F):�F$�Q#L�s/f8s&C^|�l��g ���t�"6Â��_4 �?z��h9�r~�����Y��"�&^;�i�qe;%���	�W�y*���{mٶ8p�H��o�5V1A+Z§/
c:[���#~*弖dWeW��'�|�S���JAM:��d�vŲ����h��*6�.xv4s��/u F��Ѱ�Q̚H>�ig:��f��LQ��|Δl0��) �i�O�{�V���sX�7����4rS�^�QrQ[��>
����(�G�y�ka8��'�"�|����(��S���
~Lv,�L�ZJ��,-��"���cS��L�ebGmc���� ��*�Ze�E���RVW>2��7K��9�{K�I3EY4���,�[�V��7-�\���>���0��h W�Iq1��C֝8e]}͇ԡ���xAWl����K�j�|��m�#/�m6N�B�^&T�JB�[�/��I��d��uI{^pe�)�L3�0(��������)��;�J�T�<���%z%�b�;Kw�M���rUT8;u�j����r��M�{H4$_`j����c���/K�x�lby�ij�����A0Γ����^$Q�����:0�MTF3)