// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RMnwB91DMqBgvJJ2So1aC8s6QFnma42xtnYuodvYHF72gsUTFx2tcgzN9fhchhXw
/pEc8nymtNCGYZgtsVF8idwTe7c7PPZhptqI7Q1Ay3m35GMyCa25ek+KfkGTgTCQ
7vw2Hgbg4u0QjTMbjJAPt2lKPKW9XpssfGQnEuDCT+U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21248)
Iaex3VpedulSPxJwfdH0gfOUZXUbDACOGjBU5qUOQb+5enjAa+/EUKGk3dGG3Jqp
iS0d0FkiiBnsG4gf6EprTSyEPE74ij5lu+toql19z58jHsRX8oTaEmdwesGZ4EDN
4HslJ0gKwYxRMYTK9fmNFkVu3Q4lZCYiFnF8TNEjlBtEyOgjrMMI1AnS/p6M+7yL
PdsEplHxuP0cE+KQYR6b3Tohg7KMqxPq0IUTkFg1GgOQoAnohUGdcnl9U5DFKO7J
tKPoFW08odewO30EqhQC4OkTMexw55spMnyHHspr4dJQqkcK2WF0mM/lB3voyiwO
jDqttzWsmP8incxiNt3qY84Wv05APlEZvw8uPS9Eyise4kAjQJjjyBLVWNfoNmZc
290/JqdssMo1cpN5kuRBWrVtw6tbUSjGjAJ3dU6GZpUpl7AzXiYCaWMyGGD7458X
tVnYAtKFUcgeOTqT6kDjTKKWuHGdyFMnKEuQeF0Q9CqOI7SxHfURIndsyPyC8kGY
4o/+Pf3vqNi1aKI6jIpp+P/uhSV2l06VGMsCXTF+RD9T1utoTt+7Z6LbDDItB2JU
2lVxI3Vl2/wJcZcXGzJT4CJVYs/5XaikbnMlaN3wSHCBvmRTnJ7brDrZxzd5C+Gn
6Z91uYPk1yNq/gmfjAm0NBOvAlY4aSho1K85HoLlVPlPH2jrfhIlWBggp8zbQ/0c
nkPs3quWz8sc50YxIHP86RbRTzK32ZXRBhcB28+1+gpU7vgDxpnuvXor+Jl5vl9N
IkoE3RDCGDhLIuPPBxKDlEceDwOT0TU2HAjh9ZsUuQ5wVVtKkmc0QdFiK2+fMMVX
BZNqKTxO/JihgJxwpcIt3G8BC4aiygm1cJ9AQu+y/tDbJxbIo/JGOyZ0kxKsq1kM
Q9ncTAJDNkaDDMiSKbU61u0Nq9rJKTf5k3kMHQg4Ec1EfQavG+tm61GiHOB1nBFh
6/aqCYnhfQ5VsKR3JpmEL2jbxRCTNe0h+bAY82kTSS4dmvytoPa5i/ZDEntcpsHk
ZwOr+6AdOcxyIjMGaz73ri1Ukdl7notjKHP1O6IN3X0WJvogbwlidAuJTCwTkEAN
r/zHZE2N2mwWsFtnWMLWqQTbJmjPwkT+v4ie9TWGpw2e7FvLD92GAYorLyalSJKG
6s0SoO2Wwz+g3hvPQvhIw37p3tXi5eNkqOY/mMEsudTejC1v6WjLp2ZlS7FTutuS
1PMdMoK+GxlyHVXnqD5vWkw+cPLrMAden2DX3ryAIvsGALH5QycAk/tfSy3gAXQf
tVndOIpriB7oeigWuMcYZJzFAXYYktRHrGfT4h7yUKb2c8CcLhaN6mYJiCA6Qkhy
GEaLVb/mwSB1Ok7qkUUTnigW7GAoxG+ISrnwMe30BlOma6bAG25I+R5n+eupdVPN
p3YBnyrcNiKQKz23mzccJYSwxU2Hyfdm7GxXd80vJvVUTHmwTgXaow3y9NO0898B
HcI8vI+wjKAwADw9E9sf/B5Pa0dxy36icJcWDG96bT5T3wzxWHLRZMNeiNTwv1q9
PRyzPzZr0tL7CI88I7LEESNJ9tS0vHBaYpWpfLcHcKBlKeA0WsJShYjMFx8AjIve
GRLCnXmXT6Fq/FfMhJz4pYUigd+iONRU/PiqK2NheFCymoM8xw+cL0C8w1PTccXD
AfJoQHm5IwGTmSepqzb9vU9GWwk2DiDmW7Jb6eX8XuV3NA/XSiTV71T1EAQeuC4P
EzSLJeZCSSE+RjO1PQPnVaTZ5jpyMJxp9WEXD2ddtnvS/Ntuj/wVfOvbtqGLRVv1
4GQDmJW0/1NYObkkYqWz7RkG3wgz6lp9u6gp3hUv5tqzWSqhNfaWgkwwfWsbgFA3
gcb6naM6BzOvJGJIoX17FpksKPQfILIK4/J49V0bkQTHU/JJGpN2BcQ2/1Yo1QJp
vVEOUqg15b2bhE3nLaficmKBZkTIp9OPa47ezDJ6BgcLSHo3LZ9RTbZzxcp/XRDK
WdcFXdhyJ+weFTzck8f7v4WTnwMxK8gn2jKF8pvpCF2jvnsvJ/qiepnFrtjDrUA5
7vWk5IaKR1Ty/dQXmTTYLUipQTUy+iquigmj6LORYC4OvBdZLu9Szn0VXZbBSvsO
EeV7T1NyPSEGGKiCsJJZrDik+LIZck9ryOpej2rvbbB0NQmKhsj9wDCzQqnQXd/m
Zve8a9lIQWUWmP0HBAdBFREs6ug7U4DobBu5qklwXIDzrXbcGm6KX9KigPeICDlq
gwE979Goap2dnP9AZauhkLFrwY9EFR0y6aXK7Wn3TCIf6NLX25xO/mscvj0r+Quu
Bf1iRDTTqN3lnqk6dd2Bon6QXwxeQt6ah1Ihh4E/JHrfD9t6RAxlOx/80jgXAkxn
PWbgDI3/axRv3kJW4fmDgFnURugbbh+W0wTRvsK93SSCqbjcow9FWhfE/fpIczco
zXdJ604PcRxe5yGhaWvRmP6zkrNWbxUk/+pDJUk15CZ0mVNzzDvKaJPY64AVUdjF
E/iOA7qYso3lCg8ImEkqMZ/ngtFreIP7o7xjr1XxErMF5jpYD4PcJrfnchDY3X/S
ZCOO9RGMuHV8yKsHtEgJV7nNSOtqJtHyzvkzUpbEvV0lMRD+OdHIDPRG33L6QLk0
/7co7P/gCowt/P2iLrc3fD10sbmG9ZyYqHWa4c6jgqyo5a+x0ILndd5pOIBzz9wA
g2TJgJZssqdj8PqkN+Dn/74sceTsN4swhSCpJKwJXNzFsSUe4wuBBTBjPciLRvNB
BGYe3MbPlM6Wr/FWuh8ilzDwdYiYl6QO0qfH3/Pt/AvWlPkVfgityoJc1mL2Ltzi
4q9o4sjAN+5i9zZf1QuYIIfrcuhUfxMsCrmlS5fw64UesYRlYTFJytDaZaxSNKxW
heoNCYoF0x2X7QBwtF/76Hxz6zl+MBZnELZKsqvhim1mryleu0MrGYX84pIUb3iq
x+uQLtkWpzcflo/awPQ6RvVruvfpHSCozZYwYc0n2ESG5M2Bv7q9mkRq/wPrsjGK
My1Fe4sVTYWLGEJGLvfVuQc97dTS9s/R/amHQyG/Cok1QxwzXTgoGfj18dSIWgX3
JbU/sB6xlWgLP+l/Wls6eXwxl3BC9mBnBcGwN5X0w35dJbwWQvo/epN3nBwjEnc/
sEgE8okgYdxxqrXtUdLEJNOutUF4gPLsufYzrVGtr0TWptSYR7CbXfwmCkHK8KH4
F71kohA+QsnMxvTqrth4F37eHrsu64BIX+rK+PbyXAU2ggQdJwNiU7CR6DEqOzxg
RG3oXvKSJRMGqos2dFl5v9f3hW0yp2woP+TOVAPOnTRvobgsdC6Rd669yoSm4kWl
rrVf1bEO+A59OSJmhCjaesfZQXz5Q3kgb7UW8R1Xr4JvZlatcBVaq+pRubk7lrRg
vLSX2LFQR8xihjRr5Oay9z+fOh3Uf6suhlSZqsTZOI+SJ6dca5T3L6gtAjYBm8ry
aBPrEUE8e7zU+vP7/Ff9ksL6SSkIoHswD31Y6R1erQSGwCa/o0zI+IjUon/QvlAk
7XN1EHPm2GXG1sz8CGA8j+ac8yghVOSFdgPlxn6izbp0PynT7bnXrvhnvi/ZkV5A
uNwf5YHhVyOCSgUFI+4qob2SC4ziFAPkViU4zBSloLwzdGRGpJLFv7EH1L9Txuln
VagzoQaw+ooluSUhXkH/IqPaDrigQFWPuVAZogvf708FpjHTOa2QAawmO3ZaY1xW
2qQ1NDtH3Ftj9DbqP1KPxjD6dMP2XSuSjgIgZZBwgnSdtGPgLQN9UGKP4EjcJhVr
lgxGt7aeciedKPJbrrbCHN18ieE3agc/oaDHUYgNGegTFk8W3DQP1634yPwdSRSG
n/nToSY5rYuMPsapFw82k787BnI1NBW/OtEURiY3D0Lq7V5SKTLcKXeHgyvrWpyO
AnM+4DtNgZ/b2BdWVXmMLOZNS8WEa8E+85UZtM/ES6LIsSqMnc83w5g/kMLFF4HM
c6YzoWbOXmWXNx/LUpWhXjtyQLdJE+9CxTlgkC/GeHy4RApJE87V+uqhTqucFcSD
T55vE3knmhQTE/5r2PgPLh2Md/uNa7bYBXNr86cyusA3V10m5kGk0RaHnARPfNZR
ei1BlrlitwHYaahQ2kQkOzgJO0Kor7oAk/5eFZnUBCFbXk2z5APP3GLzHRVcTMxr
fdTI1a9El+qWm5WONdi8juR3SMtuoVOK7WeBYi45tBzuZUCgk7/jfwIrogdbV47/
C3yrtvvsxvQwW7NKBb+zn6Tnm4HHX6mXd8ZOVns56rgyndy6zqw3wU78meqM4cKI
ThfROV6d4FKVMzpArFCFyCbQZLKGi5jGZAheVm2XwMXL5No8Kb8200G4CRz9PpsN
4lfo8WYgKH+YlEeSx2l/uxeO2qswnhS5axGPdFpito36hZWn7F67rQ4cb5wEPQAR
FHtNgXxUcUOkB8Suc0/EQ+YDumO1916XSvGqVaqwuJD/oq1TzvUbPxFOdtzIr4cu
2PIrrPt0iD6Gps/VVucWxB5duxpAffer/JZtCuWbbPZfn2Nz7KxBcw21+AqgaHr+
P3xE+PHRVuFyi78W1Tty68osDFOre9EwoVnTM7D+6g2YGcD6DMrWc8K8rf7rRb+0
6zuG8enLK10ugHGq/sOPxw3kyhpATPvvw5GyasNB3YFyZtcrRhKHg83qurZab1lo
Qg0gmj2szp6tyLlpZ5uAH8gmz11q3wMbVC1OYALIcu+pccDL5ZVvaDxz5OvHFMaI
360B2WToOEs0sjePXEA3RiekNCv8a3yejxrzDXiEIBeEPPrbHVFZchSCQIUscefW
UTRMDQT4L2cCrpvOqe0qRIMk0EnjgjUnqnnHFxWBMxL6mnSirsM5OsMr/9F5nz9w
lVgcnU/HAa3/K83VY8+6a2GVVUi4Sz920w0AJkPcxb95X2nWLE3Vhf9++ttHlCZg
FDAi7dsgwHJ3ud6MQDVKf+4/Lm1roWzELAkbvtQrJA1iZDU9d7OVQBBI9IFo8FGl
JS7y8a0FBw2ybPDhQIWuuPKMSr6fCqwAdhrU+swPlpKMBzz/PkvshQQ4oM+BGCqT
ii4Vl9U7lQg6KxxaniAXfPQ+BtHlQ95uJ51Q3vSecVIUh+1cr2HmbXh/nnPhl4pD
k4GdrwABfd47vQcK0em1u/sc/tTQzJKv1nhH7A+OVLtsmiG5X+F05bmTlYNvidDe
AlXGmyhvSp85EendEdpV/mTcAN7YxYx/geJPrr8VUMA9f05qGnjtf89NGoiTXQ/B
6E4ICh9C2+pqGxYtj2WMBA5bXTWcBe8ton7H+j5l9faQyOK+g96dSUdYp7F+DV8h
tHYRr+2BhuP/0EtjTVUDZTYvNcGenfa9XT+mjshLgvpJCkSy469h5GwxEoo+m66a
L1fTwR4ngTCg1qCdg7tHudp+y/hwbjs+Fqd7N8zRdQeMX7fNw69EyaGzvZVr2FOg
fEhyJ+SN5CFgHtuMqCiQziG9C0BgPxSCEr7+LKd4h3Fg3ejFxBaStB9QzlMZZpJe
+9ReLqL+8CXxVvXA02tAqAhdCp+vs1ZkgCe5Lma+JYOXvm7whCoOu97rv6WzcSfz
WJwHqT9v3CHAh4VaaFygTX/6kC3utFTP3KpAgd21O/JXOrUx2zcn6Z1vRFPy39Ui
8Pm2ISQ6tGsz0AQKjd6D6p3yA0/5WlaR9O1+LfxIm3HMeccAiujYCX8453VamBw5
EM7CpwowdDAZC4hmo0Vf74Gs2/PEahLfEN802m3xW1sHSAZufxXfMFwIGX2p2hEz
ZOCxxYholiww4+5tzrx2UYHhi+sItHWLHuXHpK2Eud4aQCWrUPDRQdk6AE+RxztB
9yTl5RD6Ud5qWM7FrCOF4Vcbg11naqkSi8sfVDiftMQFDIbLucYIEH0qEYIxFwqw
WbNEOACd8SAFR62DhzEY1VrnLtlM2KPYK+oQREosntu/iSUnwbAw4Udxt0AD+P1y
4sLi9S93f75LxJI6VML8frDbl6d6lhtSQKFlNmuo5IlbnUuAVGs6bJ6AafUAPrcw
QTexBqzu21GVjABz9sw13OMjyuEM9UqLHyBDxuOenPpa+myCUOi/X2LSI2/ymhGf
nO+59Dlwmni3RBd8WldkZ9m0TomOGOqodKtLKwq3tDOn3VAZC4XOhvBWfVBBngdg
eeQqsMRKVUOjcAqg4MbWL9cQWsypMVFsHOg3FfdE1HuGrsgJkICC4ZqFH+KJq98h
3TQlah70P4QZSoVBlS25q8TSl3Q2IVqX8KEk9CFRAJWfT6Hz+VfAmxEICMwgQwYR
vHXJUk/AI5XzOl37qPWwtNhHcWC6l988d+7aVZEtkYLllTE0YTaVwMtN+SJAj03N
17CSEMr7zNR22SNHJmxLEtPKcIDLJxkxpZKpcBmVmZyTFGO27I720YQMMky7QYVD
rifFKjdj1o9bv0mIo69V0rH0ujSJ6EqG7NpW0Yaz3cGwd61Hq+ku1Xz8zuCNpDIi
vwq+ObwZaRhpe8boKK2g3qyYfDdCaT6ML29avzdlREjeiRMd5pJjRqy9nN0tGAM7
l76JMwZDSeKWGVo2ybsQyEuRMIT5UHNp3fPfpKgroayGRWFOJCzD3Hyr/LFgm9RS
mtxqH8WIr61UQSi1/58EyhxQh9pnOuLYhlnr3x3rn6mvpk0Qd3VmTY1D/ulduLtI
y+poNjD8WCWGMX0FXBJSPJYO+ItBW4y6CVOhxcEr43rGF3YDs3OI+vyQc6D53KR9
tzuDSvKh8/MzNVmPBcbrU9hii+aEHpSenl8b51uGESWfkDAlweUrppxq7E1+l6zA
4AtZsdVflypZ4F1J/FKWEuqhJBGnA4Jxh0EoTBBFTXKrg7n2jn0vfSLq8DA3LVUb
TVs2/TAGbnl5zewUtvwYr1/2XjZEVWjYHNP2zC5EZ6AQBvetu70cuxc0TA3QeH2x
cmfjBz50fpSAPPwbeSzqSK44SsyEN/+NESUME7umcJp9LTzzpveBL6D+l9gHOJo1
hDwy9aw1yUCecuBidpiw3Jud2T4AJLdN01r8m6+OD0IovUpUgTCd1xN5FrRr6DWo
oD9rweAThm8H8GymgzgSpQsxFb+iH+wBXaztPCnNB9eroxxy7ptoV/nDvckphBV+
rVo5P7j7Xopc82fndXwWCJ1g4GuD1m6HoFXbi2Bo9zlK4Ne/marWpmMVrCgRMdxF
hLHyRdQexSTwVehgS6AAtQeYaZDbJ8hkuKH0cyJl4jsL3w/zzECT2CpGLVju1S25
2UShBgSt4uUrAnPOtZ6uv4IZ2T777FbgPhySqN4Wk35Lv8y9i6NPf4/EGpV7IpuL
2hGI9QsMzQrmh+rafqNB7q0UZHWeh99zCcol1r5lbyk89US9OsdwWCzP91ZEgdje
efncsMSra5HCkkiUC1ZY6cGgrFBS/xZNMYzcqqVvrrmfFRwXBLpezf0z6bCKcFA7
T5MMqxJ7lT9azKdgjh57jNP9sgd1shxW/kPmifqiTQDDK5otEL8Cz7RIV8+zeBRc
tvLwsMICA6pGc0C/4j2zJES8nxf290Akzdn7S5O5b9U58As/5YXD0exO0NOcflD4
wMrEVOulEzL0nF6NnIm7VrNXwXYYr70V3kgFJGioE11xm746B9gFB8egrbW+BlCo
xgXJgV2FVqcDFKw2IiTVjGUdTN7ibXuJvHgO5RCS8FSw2ExKjjOK2voxBNak79on
8J0bXSjrBBYsDmXMVv+48cYqyCUnEu4cFgAQWC+FUvLi+NN9QNvXJISYlIofjAKX
VBrR4e0GazZZ9ar18z67yiEQSamVZPX6t+JkYAyYnvVBljGxLZvu/Z10zPoieaVO
PM2lrG0Ihn6X+BME+DliZZjji2G6qi4y1AzXVMqHKrHO9EBOqxEDslG26PrIHIg1
ccS5dUhOsNxgQQ1+Z27GbdOj0Y2+bEi2PscinfaQgp1ZE4LNM0FO6ZAx470HDCrG
cj2V3y4pPJCt0Xf2mp9gCaERJd+7szLjJWTzKNGUVJTwVw8Fy3ikOzhOt5MFtIeo
UckgPW0/y1W3bBVXGzC6wtqkeRoqUL1KjHm2OM6/bShIRgvi3qVegOBrGKDVXHNe
9gXaD26AWHzyyyHHCyMDJPLr9i36Gt1Qj+5Ddvwqzd9fVNwyRkJxqFIxdSehUThs
f8l5AxGvoWzJGx8wyY+mQSC83CZN9P721JM4ZezyknD9llqyYJSQWOfws5zgTLCs
LiWiXzyB1tUqHqDBXw4fwikmwLql3xn6+RxeE+ciUjt3VwqYQUksygbZN5iAomQp
1E9XXZC+6q1/474hhPYUHlR7O/itj6LfFnmqQYpvWXXYMpzDg4WUCc7FdFOcYTXO
lqBM+m281gYAoP+LFLnDswsjz+IYubW237EMpbdE+0jOkxSSzk/EveN7Wrbr7SiE
oiyVZOEdLTmJ01uye4AWxBGoB8wsOkxe7FK2y1cn1bOSgqdtKOlUpdZERVl12mHZ
GNk0rEDxG+M9Rr+iAdU4Fi2wd9kw6qUqaPh/+7gBNrgNruxEVH0+HG0AREMcc1FW
ro/luch+ELcRKBmFdZJgX49aW5RN3hLVkfSGAlgCfqNRMxan7vPIiq6YZZjp1mmc
2hNHVHZkYi9qhB8Gwp4IqUKItVNyxJZlzqFbmZigNCV2Pjo+6DRc2ukh7UoSlTTQ
ICCe532ECCh6VWzZ5Dwcq+b/05ph8NsCSQMQsD5QgrZlGPJNd3A1zXeGjB9hl3xm
tQXkeKbcJbCcAFfDiIz2+2Y9bQXNqskEpdzPKColTClZLX4cSLkAKoi9FD5ZI+r6
TIWngaXMLU440VxqtCKEy2lQPnLja4RUSPe4mfUU4QR+dboWI8uCPhfqCMnlY0k0
ENwv7FYnC0yFKdO9ItimNxtL68RNBoQrgDOndFuIRS6DCnIaHFVtzX/B+TMS3gQH
RgvTdG46Vcvoy/8/fl9lu320q4wVgbAhwc5aDgx/QlTeoLC2vG04crsQcq/q4E8I
7OKBQz3zVeXDrSstmG7bUhqkm1bar+Mk16omE5NBY+iLuB8XvrOo3ezF/GITJsCs
7fljfmavMHpis9WCrWW4a/Fo9RMSRHCc/EuTP1Ux9360tXNaDIypKZL7PcoQ89BT
DiyvKXUGsbwL3da1Wn8DyKUqgJOdR1vsB2Yp6oWPXKSdKqzDwRMCbhI1QNenBJb7
h6yh4Oj6J5YO3xRzUjJ330RR5omquJMCusSx6KicLGJosR4+tmxBwDHs9g8NbAzj
bQlQuR/aJ9mgCxyWS0YWFJoeY6r4DOJ0LyLsc4uE3oya9juPLgoANqvYZZcBSmJy
F54TgdtET6qPjQ98n5Ud71DCY83/tAFWzYVJq2/CVEzb5q9IGjcHXXCVgheXJgh+
Wg9SSyVKm4U/qHdk/P2ZtnrG8QMZnOi+HxRF//wr42EgoVrtjmcdFmdu1wxcR0tN
6s382CGD0/LiHTpAIYuDdJSjneJUDJxx3ZhJK4WuxBbRUGF0NnOkk3LPYNoVPlGR
AL/6zMzXkPkB1CYSj8Qdd+iRPU8pinuo2iMnJI6xsZ0hjrTd0ROocT+ERsc0+4CG
BNeMHKUKKy7ZLNKmLDb3iM5mqvXobvqb3lKxb8CiMX/N8YXP+ZmbvffZo5LEEOw3
MAh14OL5TH9RA7a1qI2LYQTSO+q0XWA9JfBeI1M0/kTtDl6pS0mNEQ+Dplx5LTsY
++5JnzguhWpfpO/tv09AWGE+XzyKqK3gQ51jDWw+ytqENismVlhG6LakYNVrO6Oj
UXiLL0C3OTY2+T1VezOQbEI17iDx36WX39xnZmaM5ahxOMFJJbxHox/QzRi6VxFi
36jNUbjr+kRXkJzLKcQ8bs5dXN5EVgMdHbPt27SNGcMu83uPdf4ksEjvj5R2h/yt
qnSGYt6Sa+7HAp14z5830lSmSZ4pi8cgSQYi0LryNY5vKrSt78BDoA1n+45BbOk4
p3L5n4aidxlm4k1ajTV1+9RoxwpMM+ahEwfKSJfSjMuwDALUUYaIuKZn1QZB1Il+
pa5AZRJiGlu+1S9R+6DUPSU5yOsCocSE5de+b/NvdCy7OSRcnrn4bVa/2iQgp1q4
b8Fxl+H0JCjFAjlTJ9UA6IxTS05W7prEVMsD2EhZUuWqb0MDSiXSUQ3Tvwwm+7XG
mJtCiOzeM3XgAwdmtN17YNIv3TnGvryMTs/hVOSy3L/lFq2N12NnX5djiWl/KRLJ
uPZC0tXlCucz7phAaz4OdySLaTVRDz3YZ8yAVSXgfXa+N1cjKyYwo4A8mrEyaSbD
PeXHy7pCGFv05FbMHSUQPxteLvB8rvlD2u5Szhj+Rf/HwgmFf5J2v+ZWSRQawVCa
PvZnKaVoW6lMfjbKE1Lj08I/KlSCooVfH5MkvcLEwyw9DnU16VDz5+PV4IfDAvRv
ERkPpCK8txtFH39R9ZmACoUtuCbCu6WAz0NfxftMwIRWNTplw8caALa1xFQtvJrQ
oOkf/ORmdyK/7s8PBIE1YPpsy6614WNP1mStvchZpaJ+awkqRINwC1gr/lLd9ngb
mi0hyvn4zJLT2//g7T2N2uehEnGX7F4Svp2G1jUe33ytzqbFLCITJ0zRjmbp/SSH
zmRDquPSES8hmsZEKM5qbxJi3JTDmRnZyqV3mtJjHMv8UVe57W8kasaKziFhM6ot
c6XqXcB2X0s4cPdWHcDqOmXnhuRATZGrXciCDwlPzgi4y+OE20iInSxn7JgsmMcM
DqH6OqU8w6XWruyuN29XR9769XH1WyAKgGXfZpDPx5lohag7cD6iZ/BRjoRM8mxU
s2mli2UmDwlgjQkAd27a9ZlsFqRZwDaO5Ky2z5f3I0Zbi5uO20Qi/9+RZjDL5Olu
HLQp02rE9yAsFlEbtGYzRuPZxLrahGRtc4QJCmDHVSzB5INwL3Hia4r0pooYlEKq
8m/CIjoHA4NFYOYDzkbGiylG10fgQwa51CowHmrwuqBrK5jXQUMe9HZ1kNpDPWA9
WvEef1cDeP8C+9YoNF7b6Ey5YmpdX0zJyMm2SeboVmbbvMmFHpQpAHJ12bMPS7Rm
gf5O3O5kOswk+bvEiKRZ41QLvcHNajVtuJ1J3g9uXBTMfwgjH6nOSQxI6wpWpo6U
8deF3RlCFdMPpt/Fp3OkkBlMtwKui2ESD5pjqHYdDordsEc9kvoulnhIqDR9+vgq
Un+vZCWh1Unm0XKcdVvvGAcQD5t01oUcKrjoyfHIVLrILDTDbxXvuweTwrqDgA8d
FlM5/RBTeKYzCip+nt8hB10LmLLWEUMFSIp9rwNa/h9Htt6VfQYYw041a+wUs/eI
jmXrv0MBBoVRVuo5grT4wHgLJlEEDRejaojpoZpIF/j5DyAusDELT9DwVudyS4cx
dIsm24zzQBZcDR/XHvFqVbD57J0vxCDYDwWOgtRGIFWuANbX23RFPkwNrkVKgccA
o26WRU6I5zfpFQbedemn7VQSSM+ZOzH77bs/N73fdlRFrPFkep4nIvJuLwCwLtqa
Ae7JtOANnzb4YpTo3+fnP2d0ZOh8yBWcaagD/utaP1138oYkpUUY56sn8XZcGp0I
RCo+2DDnGMPLkhSaom6RJENV+T0SBPdR3ZB1pen7zH9oy98ixILC0reP5KTKjzsu
mQ1TiWvdzNQYwuBEGqlQEgODEKRKn5TEDexsrnx931zjWLydWNXlC3y9s5Sq/j9t
Rv7mHmxL0b6tOPCKkbws0iAdj1amz/iK31qdAXr5N1DvyQg8BInvdpGNK0Px0NW0
PHdd3dntrvKWhozf2S8Bfrj4ZUnhe2b7tNIYvf5plH3Mo63LF3e5rwHIsi9Dyj7B
nwmzG7cccphUe8RjUco/qCFCqU1NyX8dF5dEre5UFRUfC9GS8nLYLzOW+srcrNPG
kkQ3VWzMNK90MgOokyQLoB28neB0zpHZ+XK8ZrTJLxYNoV2Od4LYXnPtSB/R29aJ
LVOQurwBwEmKWYEWu5Yh3lvO1gSvvajV/n5CekpmwOfKWEGFOOqinAVwvlXPP/91
QtZlmc4u1ZnfNiTJvxK3ODQA51gBkscrYkJtxlA4C6MI6lnWw1braciAgP4id7v+
+y5WTWkcxbbTBB58OEfy9oCzVJRYB8wy+gAmhxdyPCRbDT7S9p/oPAzIMOXSnQ+W
JDlNG48lP5I9gTRvTVT1XIDG4U8f4qzJT91RtXmlVMhTiMAQn5H48yzzc5Jte7LD
ZtD4DtPwPX/+bPsRQp2UJAKDKMd0CFGujbo6mP7fNfx/ANEgLR2SqlVBTy2ePNBe
43Rnh2uOPvusKzaDy4oXE6rJd50LURR7GxduRSJfKWSbLX3Fx9P6N9jvAxp/QrT/
Rbc1VNornYay8I04Cqyzom5b2+eNJrGxGkXP75cu+RoTFRMbDdSakCrFJuI+b+nI
GosIzr8nTZ0ahIHhai6DmfOXhNjQF59tiQO5nNRF1I/F1iuj6/72u7PxfU0xl3mE
IrObuPzw5mgnXyedrqGw87tOGySfdefBvRtYMV2JQ26upQVLgfyllyaPm4MnBmKL
h7SnGLIrwY5pMAZSc82B+WGSMWFyJD6NdVFsQhJx35+f0jq52xbFK/aWaHq8wBUj
8iHDXJA1WlZQ2xECpPgaCgNESsoq0VT1+NfFwWmJAFZmYSxuFIgIPJVAbdvA+B2+
bYkQfrmE8BLUGKvLjmG1kGB8KuyZNazfGegDQ2dKXciVrCS8x7uoKZzkAkXbZbnM
CPrxKpvgGnv4POSUsv2OrtpFKEWQIxoW5CX09vtIt/uauxV7v898fkGdQ8jmNypA
PSCD00RmooiWZYZ0m3kTVgm4JDywebt3aUSULhjbUrVkZODPWylp1Wk+9nmw4d77
jmIKIIsOul0sVKbNpXGJU032Qqg1MaHRvo+vWrILNIcdX1Ue3KgNC5Om9nk0fRbU
7uEA3muSPO+s6oXbmBsJS/UiAbMCcZx7qNI2ulp4UWFQFM35+Nf5YbadOM4Om4F8
xQHRhQABAPQi1iiZIfPsIsAxFU3LZ0pXXTX3ent587qfp1hUiFj2w3bnlnjTwSav
AhMMGtUq23KNoEsvK+gruuPC1iEk1WU9s5UNOVJcZX/LWmR0D8fApYj1KmkGLT2k
SAPtrplIpaxULJenAbIC8rShC35+USFkBTsiW4aqkyyx/TO98SIEzBcmwa+BZDnn
IhVuXlt3dommhKFh4iCaoxOCXDBf1ejQsznxCsf2OZaGTKdjuOvDtbPKTleBjqLP
vBlvDDVJbQhsRupNEAQ7yOijRCdVJKh45p/RAnbu8GP11E5zXd/tOxBjA1Panc1f
biioIVGnTYQQhilyWJX09mUxxIisU4ZfD5+EYMc9a0XkrLQdNRk7YBOVFWvzkxl8
djgtHr8+aAKHyG5Cr9EAkdBMJSs9po6E/+PzlDQBSlKePeATNKxF6IpPjmLEDVqn
8u57u/bXfb7SB76DJNtsFQ1zY8lzMlQ4t/A2eXsEmrVwLEulWBTnnvjLDznxa9ks
KQ/xyoEeo/G3owfIcKmvujTXZz3EwQKVT6soe0cOA43qU1K1c5ysFqCL/3vKHEP/
n3bsdW+WZQaqdivx+c/DKFo7ow+JGBx8JHiMNGRHY0rG9t7XWQ0zgLWn5WbB1fim
Q2h3+4VdVaXTY7q9Iw+mJmbc6SDLfPEiVyEmvmS5DskzkC4O8xGUvFnzR3Nc0hwT
jm8ab09xIeEgKgEzvSG48tQjpuVsR/H6Hm329q4yrAB9Ba9tnuyj/Tl5AN/JEKcq
wfXEzPAummc+nZu4RaMH62Pd1j2RLgPxnXvsMNqxuaLxGcYJiASbqHLXFM0Esu+b
04sWJ/C5hCT4HfKIRLpK1I/NP0opq8dj+mZSFxKUE5IuKcODDCfRx/Q4kgPT27En
sZC1IRiwm4KWEOKouzZIqnZobvyWOorpnh8Amz9HcYC9TLTDI9QMeQrYDS4Il9ZR
k5itdoTM4iaN9StuPZlSAWsgapdfe1N3OJ2l5oajBpQj6taF2sbK06v+zdH4wKju
7ikZQk9T02nmTyBjOk2e7MHBRZfgXBNdpqNcl5R5sfJPuILvhCbbPQsOCscnf6qq
DhL2xVsu0pEX9VjBOe9lhZZmZfY8SNoyqj9jx30HUSLIO7NIOnZcOXsEfBOdvhEI
C5r8b13oAHVQDwXQkXH1xed5e/1Zl/iowamEKjBVrTfhDKUDupp1P+Wrdp2Nu6zh
iShBmLfBCX8UvQA8nIBbtgyVTnaVarQ13zYl2OTNdsU34onRDKjd57QoZ8EJF29K
HRDL9f/i/5hltHotvSnXVsMYCiwRuH/e0PZSA84DK6UYh1cknfYhlvushT+TYDKf
0q2G8rf0loWy+03/TEnosMu2tu0eUjO91fcWfwunhv0ZGtv2ZfhtIH16NYPrzCF0
lMr4iDJ3BW7yUqaorhXWMzjv6pMMTGIPmsAJHV5NAUIyFb+vpD+fI6QBLQIUW9+2
VkAGlKKQOyRuILQvcUh/yOnzWWJ0wFejdIbWi3rxPnxQR9sGWXU7RKzi+jYlKn4p
JPUch3/2cnJTG5ks8n7I4RKNCsL6qqdsDWnVtYdH6On6JhMBf6jESFJjahrpEVpN
xGizfxVYG5qvYbHKYVvQt5S1153hqfHHhOdjohCPIYvoBaAkmG0cRQDJkEnkhzgx
NN/XK0ppI8FLhFd9UyFoiQ7QpKyRrniPGMyghtddPEPmRsQw7cqJQUdqDBN0IVvX
olJg097XmMkqtgIRCM7OWQfgWqJwY0GQzWjYjBFBpDJD06W0y8ODpeEObAW+lVVp
iuHkfL0O8xlU5OyvjEFkpzYrgk7leiwNWJSlC+PCOe0SzkO7h5zAOYZoW3W3mgnc
XW0myF6LcelS2F9ZMXqqzK/7rhl4DE//8d+aHOQDNzng2hffvhdNcDpHMdMpCOkZ
A+GolvaFLd2FD5Dq3J5wX5maeMXrWZAwtwyq0OwBsVqW613u9oZs11zxxPbJuE+t
SOu2HcICZHSgGOLamsJbDLNVohzxnpp/VlT+NnA4idJWa8bolGfb8RGHG/kPuoE2
melV2iQrMBIZke8XPicNXUNYxy/FLgnswszS7dmGapP25E8aSTLVu73tkzdrHfpn
n3f2QARddEcXFRgR0hnYCZPYPpupsWEt/CZD/sNQl8uoBZ5HmYJOB4KMvIPH9BL1
cZcCTvE2vXAryNq9WY6FKNFc6E0KZrsKhvRN4KFt8zu6k/NTCCJAy5LDh541nM+8
fdaIjw8PtXsw/OgibWwVPwsiBAMDLOmBMPdpDB8IRDo0aoLVOgq62U/UC2VgF/am
OYCzp46D6hFNyxhRKov2jXkZ4bKyxIad6tjQ3FKzYJ5GokIVaFbI4WOl3fgKfyc4
B/LzOte0kR1aSrbTonfCl36eAZtJ06XUWD7WbR6ALAVTa3hvAQ0xOM2NlD0+ArC+
06jSG1AKz/oreUKLBs9XIumcyIUzogYCnAyIItp1Y1ykMJAoGWw2nEffcnzF55Gw
lVs0WiutiNGUEXyCwy/MlWdzvKhYLVOK4ahQmEvHfsi+/Hs7EGJWIvI2zWRTCVuA
PaazQJIHjH2E8lmkUel0xCDUC+yV7KQFXr5Szicc6CTcOoPwm8HMtxOWb3hgexLU
mb6JNkXGfTvoIBTdoS8KsXkX24rihTA2BAN2O/YMBpyP1EfUg/ahHSmBrL/imo+d
anNkR5QsLv/LLQLc3oWbS5dyqN1o++w3JBVyZt+Z7vhqR6mMvvAYNlouCy+sI43V
WKm4K9IfXwMzzQBci3pHsFE7UyKnHY6Xhn+BYGy5mtvKp9S5vE/LcnfF3dr+UjIm
DbD6l/7Iq1v7ffxGoyWZpNvAOqitKzjY0NKn512r2Azi3NdNDyrd47bmdK9ib0LJ
a/zjhEa3BPNNqwrDFdIJKgVb+9lbWK9PgnCIfGdtiwatkhVvtOG/a2PFNHdxrS1m
FF9xAVO22EZJY30/oqBbMQhxKvmdg0OJpWlmbJmkQQhhDv4LmB1NVSOF1LNo9vBl
Ac+7OV9jxU44APDMwQ7Ea8J30Ss0M4D76RuNntRzw7f68yJUrbX1sqA8yvy0M/88
M3OUZVvTIyAAn0dpV8qbw98Fb8XxwDnRKoWC0PHJcM22MU0C/VlotCAGnl317YDn
yVrUXKARrTUjm1ht/M3vw1Gg6cjz61wmuylmHKDCk/6pCTa6KGeMWCO7DBzm69fV
aeWFvI/S0jph7RE2Ct5nt5KRScxeH4dIAZ5Qpy5BXDcXj0e+bxhWOUsP/xvmnctP
JinjEBDXvgqxZ6b1Pn9ISHt44xk8EWu4kO5iCoKMqHjbYtPEMWyjsLsVh53aVaAQ
U/NnxFPzkFCC0YFTDzbvHRWgFwNpDvoy3RV2eApph2yr9A09nOV6sWHE6sXpEqNB
Er7RNPoYXqA5yoL7Nls0pC1vDT5ZcumBsBw6CRnN4D80FP9Q5aX9aJ5iYC/pa4HH
0yrqc9Z/LboOikFpelv3HhTI9dcsvjz386Mjpd3YNcTfitXGJ0+DLTe2diw3pElu
awnOwIdlmFCSYdg5FVlg3WbjhdhtSKAJlFwJfBAPOSvjAgj4wOKXMCcffeLEEbTc
qWoO9jF/yVonVznOyYbn7kYzzHpZzE/cIzoa9w074jhfTsmuCItzcZfrV+6Oli+q
qLr5bmpUvjVPwUi91dSd6PK4J82P/F6XCHnuzkumD93+EGm1FqLdTwxupbyXY3yq
gRuZGYpbX66ho4vKZ6A0rotFMnFTU2Z22tk20SXYlBDi0IfQ6blfqBu6yvBsJIY2
cBFl9soSQ+X2Y2SMhYA8Eio03lPjz81q7zrqKF9QfXyzo0xeguBagBDLNq7JAX5k
B8juu8rdqmVwliCEWbaadP0A0O3yg0M1BMSueNsEeJmtuVW6NDDd81KLXeRBEdqL
bb20kdB8UsSVViQUaQdUB/Sst8WIyaszeo3tf9P3Ym0wiV4lnFv91NkcLsUdg5ND
lQtLh1phzLF23mPttwQmCbyPHxCwkBOPgA4ekckiYXeDEW1q6V4pt+JrIMgdZSOe
Ky8D5ysKyT4+TRi+kr10epSHgownIjjn9AVfWc4HogCV5PzkxY9ilyHAH58HOfB+
U3ItyLs8Z1Rn47lGIII4iBrMZ4UWfEdXyCNBbbxYdnDCzbMLVhYW7UXEAbxLBJm5
iTJVk0+flS4oY84dBL5w4gds5xZKVnaRYm4mz3AmEVhS9NPiqypO4lNMEwC1b755
nSDaoaj56VwIXNVBqQ+E4N6yLqm4xSxeyqSMc/RcOD8fvLPm2hWCQdNHcLJ9e96z
h92w/5hHNstMVczzAddmuyWSgFgDJw9G46zywm4S3dLsBxBUDa2dZWHNNIcaMJ33
GaXAqkw3Dbff1fe7g0W7YKdHGs7hNbYmQ/Oy2Sx4mk2DIHvCF76CS2rk3rvlunVx
iajnt2y29UEGDUnN/RjKKRvCOVkMs9I2EKSg3P3sp37N1E6iB31UHldOl2129wKN
ZoK1caxp6JG/ucAw4eGeaIOVoT4TtVPhfn6B7mxy5b7Vn7gBf/TlgGNNLTV+lJM+
RI1cLvvQfkuM7+Hse+2657xMnUsvcd1OG0NodQ/mYlue0z7FWnWx1AqKDRwotKqq
RB6YnbaMtO3NvffmcYHuYRalAr2jqniUUm4LcqVoqKzn0ec+cmdjbGkhkj8+rDt6
BkQm9t3dwXGcaKA+aIjFbxy7FAPYeHUJU9CFaz0gDngLEjPs6ZeB4EULV+DIY4ZU
x0lgER780+Wu7dTr3428uP0Id6cg63x7BPIDvI8C1vjb4CFTv793vo7ZwkFWaeAS
VZ29bqGhRujr4Me1B16W/tpHbGLnHYuCDnY/EASxqyNMhJnhg3ZP6GuqYkfVCUbn
dz1vFUac7/SgaoJN70BSCUKVTR0TBTCu7gRR9DxCbzt95DaOjztR17nKunBtXO1p
C6W/ytUUiDkFRpCv9i9lAf0X7ZAz1ZgHi/cACqke2HJz5/r2Yo0mLuDLQteQyOjh
VUgAOJ8L75GZ6oBYRd5eBjnr+8j7TWKHoKxBx6mTd4v70W8Jni95kDhGVaG5W/ww
GI0nKF3imGx6dnHm1/j6U6TnKop0HZEpPMdnu12BW4rqZsCtPy2jdwxt74edUe+Y
hdIXPFHMNp1m1AgiBfjczXBuMVcTtAMIgqAA0iIaJwo/5zcXhbtNBPMtSeIyksN9
MPZv64aoGi+2GbrHEIGH2/RZ5+IHrVqPRSb2Aae7lZZpXNocj4btEyrXcdgMtyop
dzxrpl5Nn4hIOBE0EqH7I1VK4kpBCuXlsslzit4EHuSEfAA4rvDAOdLH/9EqQ5Wz
/nt8odyfg2ijgzb3CWrPAi+RbcBePdy00qs5IApWcKME00yk6+ou5YKbNMSX341M
hKDqcOx3iHqZTxcPK7EoKc6YpMGMUHnyD2OGjSB6ZKFGuAEKwaUnPl3MWBFgVIwz
IVRSAW+zqkE5j7kJNZ2EX3MJAaZTwMnmyIjr2ex1DsclQuEhRlMMLt0cHFiaWrfI
xqQi5OQpTnNeSWN0lATsFXlO6Yg5Td1BanJagSqywASOyZBDh7wB4QQ3qTqE/oxb
iTTslgDlxq6WwoFHA+kV4cL6HxjsnxwK/AMOikE7o+H9t3b6vozkZgOLwTaAKMXA
89Jgwqq39kjU9qoxQg/KQWz2X8qLU+uayPAz8X1L3iXemMizzBB0ACGm7c9R3tr3
qkjlMuN07WlCmozEchiVIbVcua9qKDlUy+c5Qi85o2wiKA1K3t4YRjX5wkoWCeUo
8/o5WQyTwp7CNVtHzncz9NyxfsMf5J1s1/tusaJpxXWbV4VuUFtNxDQN4OczSmNR
qukBbSGxAwbn+FLR0LqBQTWoPrUx1kSSjdsnY2YoOG7aC5Jb3c4z7YqrlPk5Rk2S
jZHpRfp9x9NZFzxCMWFVE/vLMuxKtaE7AyCqOICf9/zDpv0nmX2VEN+VBD2ALzVD
yo3+g+jbKPdxHWdm80UsXAOtIviHRvO9QQE4nj9qhDguSlb03IQJIevcXKLrbRIt
RfJisdvhpoEOPJTuPgdPsBsMuuL3/+duIWj9cqUrhqKLIfp9fjGDSPqgE8eqvJ50
adfOc1wO6c3ty1fFwILGEhvU9MxlT2F5FYhUN1H7zpTjxlj0J9ta6jLuIsMYRL3z
W4OtxYNT1W8djijK727UfFgDLsg2WMt0yX4RsPGbGaol5PW9WV1FE0bFxtXz/GFz
RcCcKT4+/KCtDjnnSI6mo82MlnR5ftzcdMnDEkNkKu4erM+VARuL4nkKGy9W9jZx
BC/C9ldfjCfI7kWunfYvG7n5GX/w9MpJOipH3L4RPhAmDULc5VTLPGdRnIsgW7Vw
c9Id9SYOoJKs9c6llxAe6dW51KdkNWFoUQyy53Umvni5RpEzKRoxXahleTIBKJqE
IgkhbRuvotTUOHiei4Nt9Ckj9j53MCuIMDoZWmW7YwVzG7sQ2sZDSDudElzqErdl
SmYwhmC/pWBl8V74Cg0SGV/8LbZ68DSujkBxdj0iui+mZcTNykkIL+W1vFHP1ldh
9YgWRvjToroZVMQRWfGb4zdN7rskAlDLo14bDSHcs+4SVl23nKpotuFcqOAf4bMy
gXcYTAxdeK4VkROQAyALJkN759Xc0no9oOyagiHAYSRg4hxyyz1nuEueHk+YdK5d
bDPqw6gJbMeV3ES6O+KIj6R0Eq8CuwJ48gDTO0ow4SlADq6GeTuEr1LlT2GcP6ph
ptoRh+qPjQCuAmJmmXVDZFqWICcKHdSo3NzJX14Odn0/Ei3SBb5JJfb7vhGYcnQq
2A0h2yYUljXSbJai1BsTaVKW+yK1FAduGbURr0/H6jTI32g7QLv+tVXepIfbTgF1
ff7phW+q9Pgn+1CnTyqFn8PwxgAFnlG0LdWGyytXulhLkTeGtKazoaJ619v+M9rQ
pPmWb3dGgYsEG/fsYsZnXEwFlELkBwLu75ZTR6S3iGXl8GtGtloYXMAqgcadomG/
/kCNN1UNzwOhCff7IU7rDeVv+5p0H5bl90XORe+0UeHrpc70jcovof3N4oqQ2Cfd
2x6mxdZFR8Nvtu6DXMcow+rfMNfNjpQMZx+OKiTQk1kYVeRYwxNMXXEoNs2Rq1I7
cqrTM+IfpyPX18rI2/U1M3jMC9Ky9kTmLae6f/pCzrogGBOYYQ6XRyVrIPq54eCX
8F1IYXNqDMqL1EvKxCkFyMATuON8YiX8K9BqRk5RF9wfoWX/4aNJ0FByDohvyapt
cfx8DtMb509PweIFL+9j6bkalllgXtCCRo1PSlbQMzTq8X6pvq0yIVUXGLp9KGnq
phjeB4wqZZM7hOBPl6t77IpC9ntBiC4lQilFeTUfnLodtp5gIjCui3NM9fN6VUHv
2jdm87+2evnJcCqkTA8KixA8PB+hHeMdk+9cYI0BMUA2gsMBwcEO4UVhXz+nu9Co
rMEJY7NE9cUOxb39uSadPMi3KsvvoNQuoSstNM1oNvR2mn3tAM6L3lJQlMtj5HCi
yssf6mXJ3BTwzuuBe+RS8nN0rIX62nlOqFwnATuJ8+kJJPGIDGwdfzDWUvcCcfwB
tqnzxibsu/YMQFRoxoNOhd2L8MuasM1wJiY/xpHfj7e9/cVV4GtqkBiPMR97pqsC
BPajfd4875verrGz5QHoX7AZ9zLw1l0pnL6MOxMkAfjYk8/mRVOdrpjBcKAgAToI
sXdaqKfetseJWb3SxF7MCEz8q66EuMv4LcSQ4cv3dzsAoH9Sfn3Sj/M4f0AVFaen
me65wbV8fEDvgtQ7rzDe2s6yxhbDDp2C5S1i7NB3DlC+r9r3laavIDm84lvsmkV4
iQ488Wgj74sFHec8H3sBa0ELDMN+k8zB1ddHC7IpGzMfR7pjgK/YmuzTUgzpAJMu
A+KHeSMbGL81CGx+T63tDNHDwb1rJCx5LW/dytfC4qx0SY5o/mU/3iI/fF9jY9q5
c8u/U8ylH3HSG2RB7iyVJ8ynlbgp0BUFQYcw7pF3qAeF7rBnFTiMWV0hq1rftQst
Y4U2l1OQWROFmpfjiTeFdiD83csz6yMJ2wW1s8A16CEce4DVxHTFFc8AS9thDlPG
m4sOlXQGsPuRaoVsSurCqa9ywGktvUGdpTGJd70Ng6o3YmNt1cwqgSXJgluLDkEd
p3E0GhQn1ElVyRRtGfyhKhscBkHGf8F9ZBQAhhwwQKu0UhEQ9o6219+I0lzdjq3t
MnWpsfbw5KZWAlNGhVvWu7B7oOMXw0stBRpPqDEz99DZj4sWbKxXN8uLOQ+xXScX
q0s5/lasVYSVEAzSko3wFd9vlr705WKxvYOrFF3wqD9v4JBHhS8nG2XneUHh+oUk
Z94iSv4nrib2bq6EObF6dFFjD3sN5iz2A9ONJupBpEioiQWOpthdrk/gN2tpcx8Z
UudVZJeSswcMXe9ruWCVe+nFNDFSYoaLAfqxNU/kRvTXX5YJgpQpvxAk/k5IBTI/
efZpO4fkkyCPBg5vZj/OQjKXVCmldGRMgUCRgdJNYtnNBFBpRRurL7lZliKAbNel
XLNyLfBwLKPMIq0or9ClFRyGTr0ZTHS0CS5qkLEGUg+YsvGgaRhUKXpqw8ndPpt4
MmsNfurltyVls2Mz/tFSrp+v8RIOrhOt8rwxZWkIxGo0o841i2rrAAoSzb0xLBw0
PVV1NxxNOK/D+rlFywdciSm5IUlfdCzY7wLW5Oo6uyHVgVuiofaoRuy4qE/xZf0Y
NTtrN/zaxcLygEtLMUAQzXNrAiEDpDpvDpQB3F0biIZ7sIoLRUfNc7lRuRsJYvMf
PHXWbrhm1MRj2y7iSkAM4GzF1uS6Q5JojH02Y97V+FhfjBSHy4r5tdafgLcw90V5
S5HiebpzdQLS9WOKQehJ1NC/8htmM6JD5UqDzOtQYpbc9hqcseDZamjWBh2PdGD8
YHJFvIMOwEiFkCZTpouNtCR8Lj+HoKItkzrXj5iL+pbstmizCpBv5+a6JhJW8hBh
oPsaDnFIWP6jR640cO2PreH//KaqOtTahU6oKtawIYgbOri1tE9qYrnHePOO+ZD7
/AhasJWbbPgKMWvQXPZD/B+nJ0zhJYpuRQkdK806pBbMSOjuy/DTPigjEQsJIoWd
+G1pzOOEYOeh7hbEoN+zbxtRDpV8SJGZVbWNGVj+z48ekhQYiLZO7V52KBgG1UcG
hyVjQZJEVpiehUEXckayBGDNoveZIvP7YVZT2+4eoz2EGtgBeaAxC0ujZUJBVCIS
LMINi876gGArMuo220Cj0SxjSS5iNDOQbcYodye6Y1UafRsmZ4zfJxy7AviCTyJe
lqZ1RqgBYcKG+5G4GSM5ko3YXpHZiTmrbbhN82Ai9TxDbWcBJxPW82pBpK50VTJf
VzXLeOS9yliveHwQduRN9vLK3LUK4nRZoicFwmjutiTSZNQ3o4VzE11rnGgKYXRq
oUSJRT92FOTWvFdxJ1wHaoJSqO3xwDwuahJV57p9mgQcRhdhIuLcIG4VT5Bg6xIB
6ZvnMZMW8K5dFX0e4XBb2g7dYeTYYnbYcN0lTGqhO3EwJsNoypdhwwZwhTtUPixm
XkveZWjQDtPrsw5o88ZmIYxWGzxEIoj8rEuN6wManu+vCYWeGKL76UR4JYOW0heS
y1TMpLFBskqFRL3PwzC7S8WYVJq1ssbcq1N7nctx5ZVud/SjREw2wbhPd3fuDv0I
a1ZzmTjOKRYYlpDHPxX4CHBw4uTRw3Z/jxapT1CtH4wKrlBO56ahh/fiqHDyWb2s
OFRLTV3UA+NJiaq0l4hViVasJDsKFQRBTYXZZOMVItBlsNtU2kQe2GESXcna8CyZ
mNJV8+mnVNL7jVn4ahyfNCo4p6EYa93NX32UklBdEajU+NtxrePX7gS6DkCQSXQt
wKFSsg+/qQ7Es7O7ZYIRYb9vwP6HnZTXKst86cdBlrMebDgNMy/tIJFpaeWPU8jT
pyWQRboXWNEbu6MEbdenrYacvgsX8QRxfx3odL693Bnc5ek9Thnb2TRYX9JtZJ6p
ZrRjy+U7NO/Hkn66ZHZrjPkpG0ZPcPMYX5cMxlSrRCxQgJyG1qkQqNLjCcIWE6aM
Nfes3F2XKTFmjfiFVoXzmcHfkRXEjJgqaU2E+Era4MK3IhkG49cq9vTQXJ8253gW
NTzsXR8UTIp2Wez2N+QotzIVwlJ7brVdSGfSNNe7v9+tDJNd7Wm5mqHq7ivy4gcN
UoAcqLSvU9//F9ZZPY/Mk1IQP0ODvgGrQdZdUMhYAym//Lbzdd7E1dILPFWy8MpH
bXG9nQA6DuJeGw06WWwLyQEdnBn8LPVJvqR5izYUsEulhHK1h+0w8ZA8YGtwyEAv
k5fPEoJklY47dLsaDIzz1ZzF9T1OPF9HLvHWEEkeQBDGf+Th317iNPse18BMAXr6
RMFNPKrvNkr9qHR+mUd94TePvqlNaRrgRtJE6O9EWWEkYo5yi5VYuWCws9z4cpmg
rwKX5ao0nVBvw6ZY9nE1J2FUzLAkumilzj72/3vnVerbg1YTINKgo2TZryIvVLSM
+VGNTwWsnVHj+4iYG/BMB5472JW6fTA6scz6w0r5dj4LmeC8QHLWVmyh615gVVzu
bo0YBKBiGVBQTR0k15HFExV/a7q6ih79dx4g8cHDLgQzt1W93I12HMpH79Z/T1G0
hBPjfIQlxR+hunt2T3tnYUnpK+rD08WTekp9yZdTCPnG+FsjAYoefanmU4tKCKK5
DvQgMldHDFtOnUarhKLAxuSlNJPTjA0DzbdVJsSHkMnQ0HeUKH6cVzfMvW2BGcS2
id6P44JWiJXZO4RP+0+p5qJsBgZ09R3LIMy5kkURLGoTtUY1vqpaV3r8A5Admv+m
Ze2/PidNtkTfBm7ChbWb7m+9f5TSgnkDoTzortMeSqmmVnBM8hB7jhcYIX+T/xXe
iT4q06+LhaGlVejgSS5rgMlXAkBO9vQg9WOyiyr3Ms/icgGqAUQ5iz+cskOW68Q2
6Q/jV4IERw1hYA40TnrxuXA0dg7n5SvlNVYIGPdDkIb7jzwYGr9NUObkIupMQ7eO
84a4/Xfyodf0CVYyMDPRYvjztvgvJytZO6eujtBcYZDw4+z9FxMu8OaNX1CzagI5
szbB+F0WylLrpS1/v+s0Aq/SV0o/KCUULYM1C44DmBwvKX1nXAt0BYcY96BkBiNc
aBlGBrrDFPUMQVzFh2Z1SzlRVizBkuninn/x683SMNOOZcVTRGKUfSqyzp9cmJC0
h84yuJT/N6XAOQTXziDx7t7XCVSmH2oqsxCrPH5X+n+s1Z+t8hkH8oMA1rixdLoC
Jjg2vtZk6pKuIN4KW846vVL+LJ1Ft9f5fpy280MiZFqi+gOgfl00pDB8etxEnw4s
Y2cuh48RFL6VJDZMj9qYJDxp7tRg5utLBJkwVHKBfaxjBCT3JFiPhhzSjYBkF2AO
CAWDUkJwAGrlfmZ4HvxLqspLC4qcNKKlOzI/+w0JmXcisR4PVu3FLaNtjmtecR0X
q2v9monxt0DfH5KVh8rQor/uvm2T7tyByn1DPw7Qen86I9Ac145oi53hWjuDzgw7
jgQ2a78JFvvu4j5PsrSxRqb8coKBIHhUltWQi/lJA5xClrKTVGLLfTVNz9lncEzy
hOPgG8i+l2TBTUHG5kAI2h6LvfSxSqW03MwdtacQ/mWpO492srYSsaMm1GESVHq1
9JGEb+o09NILdJer0CMg/7Kb+4o4XKcbyk5rWLYGiZq1/YcjEifJJHh+1v1t2FWm
ev9Y/TxH1l1DTyRAzq5LfUopbMIbhL7+Y7mnzWWvY+t1DHO9Zt1u5L9qT0yZ1kY7
UeXypj13KGXQgPf36AOQ/ZcUrKnS9azrLPV33+FCoGvgiXeVUPS+V3kZHfeLCnv/
KBIkH4coK7MLHwF2R9wTh/X+NqeaHl44bIBVsAZBzMsnM5Lq4DUlrPTKjfWwbk17
r8ENrCTnNmG63/5JXbpG2RuNAFTo6//VPFL5HkHp2PlHYiYuiB6vB/RnLCGLEoxM
TeUc51XeuDioaA34QtwgrF0BZqj0G/Ht7oK8fwvruLZWBMZYv6quVpG3haiSxbd8
VEr4A29PlhGvUunqj5+biJnCOMz0Aj7/HWAmaAM4iT1DDytQ9//dd44I1yt1Tsoz
E6CTP4mn3J4TfvkmRvtQisAzVDvEnNbKvmuEcSjHSyIWyFx9glaBnCdgPJblWeUv
EfgSPctEkCbzggEo4GkfOeRKzobHnGmMMLdc0LO5JYrrIYCNBDdOxafdZhX+5hW1
xULl9+JFTPLiunvRYPaGQRCZeleW0nRT5BHqBF3UjrS7VzR/h7KJx9u1qhV0DU/t
OG0DtLzDWHtsyjavz1tIVf0FJOn8JlefOmVQE9hORC9fAK0W7MhCQInNiy11lXFZ
m4z81QsxteTpxhwUMV6JgYMEyemjECh7WL7c0kAVkaBl5KPSrTPjB+vtZBLY/0Es
5De0VeQzeT8zYcgZXTilafeZGcpUfTsjCqjy96HQIKZb4syXDRrGLPT5dxfbZLvW
3BlbJHbKUTFR0lnqW/4rSimnxP8iF0TfzJxwfKwBEaiqh29ceZ5GndewddLXayiQ
gYCwnQdL2yAZPvpfepXsvGWUtKHRs0gQDFvwj6eld2iBDGDkoMOYHc99Y1BI8ET6
/DgBWYxTxnngbzu5aRH29nDj7nt5d9k9AbP9KodM5UVDwYIVoJZbwweGbpL6a7DB
6IxrVZNvHo9/ZSWUH8Egk23mBkx86bySBWbG1OAjd8hSO2tU3HT3tixE934aBdow
525VS2EHJbzjCH9SFKSruOdgsuOus3Qp6+MPlIMwZlDplClspCggCOGGyj8HOEM2
7gqw4rcgAEWPnMwylP66Z76tOD0s0pT76L28i5F0nkVyn/6DYNKqf5m74YQz+Zih
Li9GnOtHb53i0ZhFdQ4yrduiX2p31YMJtIMHKoi9lTmRxdaYsKi1B9Pm6SKaObID
kJz+tgPz/00lPDH4hcFFgxNzpLKpuXM8493BoPoq/7ixc1E0QKsFPIx+pa2MCvbN
y9yTa5v+qGdpqOveb3mZMJpP/u9079D45maa1+r1EsTTIFn9TCfka0/QcpVVSqv1
GLaXx6HjNm+lwA5wZZjH7M2cIyXLZeOShTCKvEgepTO3iGKRjEXvpjAELQdIW337
c0/LK6ZSn75Hx+EgiDqSzjUOZMk4AATSOxLI7Ag699YchXeNKhgtuuzg5c+lyf9a
EbPBAFey7uroyF1tPkjmYWPAjQ1fMJmaT4mz6Wo0x6xilcf/tIWBaYZFmf0OH2yQ
41YnI8NefV+2vUmlOds6BZUTbj25Hd81U/jDwDICl6SrqUhez20FTekCvuf4vOZt
wwjhFrQ8AKWOcoR6vXUr1qKhc2/N9hFr5nQtiJ7PLMzkxS1GLw68w2wA98GCB1uE
jyAw/oZKq/LFNijxiCbxoSgwaFytG0f48AuPHqOjRwCr3LE80FiDucBeKMVgpxqf
sYb67B+ZV5X0RvfQQmNvirc/+FP10Dgsns2nLeLCOR08kwxpfyqzkkxfvWJjAgxX
emsJoDPbd6GqBI+Aw6H1QsiXbHHI6v1jZ1h4AUipPOxQlX8t/9J462vzqDX3t9/b
ZF8lPaNCzGqZptPkwQrjgXJxdLWezKMQ8CcvHoqBTv3YhK+Bgf9qvf7IQVnbzHSn
S+HREaCmJIraZzxGPo3ykTE843KnJtgC9Zk00tSbvzT8nii73uhOXZ67HEuFBq/2
HaYcSvrWZ+gRdC1ESfROrHdLTi1p8Zd5MWSzqvd5GYlPYuqqxR8s6KlptarlTZO7
ovbixPI9jtojoqD1VIM6Nfmqo9CY+ECDTdGLTU/D90y4tE5TTctQlaQfreByeOca
JZ3iUiO13Y0P/fOjjkFVg+YlO/H/0SC+EDYjwqMt+bddw3an0voVmsfZf3MbfOUK
iHVLjtqyrh8NpubHHo5qxUgY+JxK263rpW7/iHrFW+59Hg6CkpnILMH1Fo+Bpnnb
ZE3Opj+cKvnZUY0bu+OpMLTD7nx4NmovhaGL+qS9lUTlo9FLV1ETwhHitF77hnCP
0cRS/zQx5ylwCXl6WUGs7Ll6pa/zD4GFqvHjRv4FsXry+vpF/0KtA7E9VarYzkDZ
RI13PAzD+xxtYgdS5GcTt44KBdBJMhEzzWAuhqs5vw/SXQZDPFLq+/aKVPuviYwh
r2hto8gfcRMsaAy+RmBEijWWBRqCNAkyZLmdCyB1e8lXlEhY8jLSB7ZIRrryRZ1K
HbxHd41dbCrBCZ/oqicTVUtLTbXxJMwIPRE9bUWUN3/npsthZMu6TDzedxbAV208
THsHpA6kWvz3f9NhfJWNt8jAXPMdoz+ysgnlCegF7T+/+lrf7K7iiAisyePLPagr
AAT3eYTlBIBq2VmYdFsfovI20IHq2p3xnhwSZxuH3MjR6l0S21Af3mn9Vcrdcs9y
ka3bNrQxjlj4k96eVx8qkgMHOOmLFAngK5AT06UKlYTPvBRySXQV3JPQXSe6LujB
2w3KZLgDLvsq6MrOYMhCfNcMCXTyugUEmZz70V7VFaKx1BrEquSmNlq9kYgFzYFY
IsOw1nrZtsYLFKbar7oam1FrfBZInfk256qpYNsCXrejjqy4OGbwGV80fE4c8KFr
3ADhCWm6GgpMbXsAFjgrPqBVUJRFdadVpY9XaiwRGtX5fTnAR5mzqiEwiVsbuB11
9Ji/s19LDyVbf6i++K+Kga6lvkwgZe+HYhmvS872vHSZ0uG3TGPbLIDpj/6qHX7A
ukrKDyl8EPfQnJQq7K+DbgOdcHSVNdGPHApBhMQThc8tlyZ102KZmEI1tiz3aBAb
v3S3eTun4wlPdtXzBiHUquseQpkNe1WFO/n67hIqG/1oboXPX7VI1C7mOj9nV+S6
rLONhqKeeDL/Dip+mT6rm9kDlC16kZQxYHW88zfbNrJ6W3PEGGBrSpNlahaDJlC6
uDRG0qQ86Co71Q1fCO3r4PkEDLPzB/0Mb9WYvd205NAPVyHRb1I1de6kaEU+Dgeo
cZj1NphGsU6MD+U9Utzvylq+MRHqt3yWFoUtnAKFLJtfBhxTJ8Y6eo/QpQEUGFo5
gOn7658uAHUhfQ2t15J37jMGiyKCb9tbwadDeDHShin3P/emsXh+RjAuWrWxONcv
CUrc+RYAOG4JT+8iicsio3ue4vWwUwS7B3Mg0KNx6GMb6SxMZiKFxMR/z+TTFiXC
C1NQRp763yAQI3zn6BBUCr/M/kWk45DQrQoOYrXzDy+UMccnsg/73kwMU9pBXHRN
xftUOButvbGgrEiHbR1u+l9GTRZ1yk2j0JV4MNaFO6nKVYZKfspG3Dk495GPRdim
FrgxD0372zMCPkgAVs+rjk/kY1s7eD2MpqbPymsoFd0FZVkvE+D/a2SkP6nuYSaN
bTCOMcWEZdQPlxvb1qUKTj9eS12q8598c9yCDzN8CsU=
`pragma protect end_protected
