// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nfyYARB7n8H0lR9R4G5vSuT8Bme+Uf56fzNgKrLt/ZV3vqfVNs5xTy0qmvhZ02A+
pg/Ef0Fc9i/xdHhifiJBuZb03HAhf6sGQ9yBclqOXPEy85e7bL6jQcDgC3vyERdO
J+Lw4TTb+QSU9mqAiNtz58tJOlWUjaD43ddbW6h3B28=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3664)
mu8KIqKjmDmbnM9YythwGECD4KmoOSel+5HgA1YHtG1Hxue6kHyIybxHP9isd5q7
yZ7mxtyHcA4mz+Cx6bqPfnoJfUJMyrZAndJedV3S7S9K1r3rDeBJFQn0jXZmndhi
rz3Hta/UMsSe/4+2AasbNWX7wdV89yjn3m90egDP+dxTrPFZJOnO5RHd2ipOVwK+
UFn3997Iuo8R6km77+wTOo1Fz5Zblx91RQPoNwhfVL5o3h8+b6haLrnxuRmw0OsD
tW3YirAHnxyuelbf2pqfCu5q2+oDITEbT32IRgtu5QDLF3EjGZ//9UTQ+R6eFEOt
+AnethSMsRxqT3Q1RmTNHYRtQhJgjiTvNPf/KY2F8Eaox0vDb+CRY42IV/V6yxcY
zNsbCW1h9g3ydoVQPelhSKN5GlntsCED0xNdn1zIMSU+gZIsqHJeudVIH8vwo0Cr
EO7j3pIlUIYNUNbO2kBWTcFKsHXHS+HXX3wmCEMx5n27GDbC22oLegI/kbHAlZvM
e78kLXEYUfEXqAp+N5zkkxLobwiFCHXoJHDvY9XsTXjzRyAkb7TehTr828oqTML9
5GAaEpsz6XA3VGTvse/pwIUnTKOvMX8RKtjSFxhAsFN+WumObdXbcPh2oZw5SW/k
tGXxPqSWOLVsvJWCP5hjpRtVSqdHHfcr5W9UGB4ID6xMSROBPb1pW4ICWNndo9Ya
M8PpScrB17lqhsGaKrxGICmUJDdBLo7Xl0SqRl9pD5XmeL4bZmyukBG9cnsI3Tel
ujbcGMRvPh7YQB9cMearciyLAuwzqdH0HeYkj4eRd9plIwnLXoE9lJXo+G2v+4n3
SKPdmiMyUi6Yp3UXDBuA1O20G/qmAlkm/kTwGBhtEp61v1BXpWBM5pqm53AyoqWi
WI9DIPOBClbCNuvPHIY4YAXbVOzy1MrJZndefrbK6b8WCl2DufMUbo9wrASgOTLo
d9Ra/uQNHaAzuejSJcZ4QiPhXZLTYZ2OWLSKcZX+X2jI0fKWhuFq6Wh6doRn3ffE
I176LB+v9lmhZMNYmmvuqx6vKs/2BQXC/R63CxynRmabCmTV/YQEknSvwFX7AI74
xmUtZ3/fQIweAAZ6SMAsuI+TgMtrYJ4ercK6vSyCiKHovazhD22VIpzdLnKVrv88
uQgcZCim2KsEoMS40DIih/I0iQ9rpboLX84o1Hc1jBd+WS8sBYe37YDfwy2vAd+j
637UA68fj8YCu2MNlHEj7ahTppT/P/RgJ+76D4yfm2zZurhJ1rFUVxp0buEavjsy
yx8C5oeQpuftBL4obmHFnnLqDv7MT6LtwkZOmv5Wvvx7djo5JDghPg5LSe0DPzUL
bav6tnMpWx/yNxyXhznG8/QGUPIQdiHZWDxOIfkhyB6ZtQhY4P4os83ENUX+W/EK
jiZVb2vV4mAvdyy/YnE5s+Xju9oqzLWYjrYicGBqIu9NbCnjduCBClwZt+llabjn
dlG8ggcqtN+84a6HGfcEALRh1dxAhXL1pC1oWw0dN2n6FhIbsYQnxW8ns+NbWasU
GeLXJsb9vnh/Zc3KR/Gd6yUtSQemR7jWyQbn6cG3MbrdiXVvYu3Oyn1j0CXUX8CY
f0BzX3RsIutpxX8KFV9RXdZ6Zsqh1yTme5ul1EhuV6jxIw/9BTaP6hVBQdJfJvRo
zVJhp8qIAovSmrKVVY3g6hBmCnpgd4047U6kHfHQcq9DncB5UArhS5eXAJEAs3uz
iymt+url5TMG8unGa9GqOLUCYk2huF3sEKYuw495ZsQov1Lsjz+WVZfjAX2pgs2A
700sSSi49P3aay3cgohZe9SXKLo6b/1ogJv8NOXdzcZWCo4Eg55AFW5GImgs3R7B
+jgisSdd6W/ffbfwjYrE5DkIMEVOeiWkZjcAc+hxFUghOQ47jJ7CfMmInGU4LZ0J
gxKEaL0n/vyGQI+P276y+niSeFelwQ7NBth55l2OmgbsP79nPAVRyhLXd4p/u3QP
m9E8w0m0TGw7LfKxrZosbaXzJjKIFhgdZuDQHqcjBoOzGxawBnKcRFa2+hwGrIn0
I2B/c7HsJExWVGdqXWNyCqqEklXR8Ci0IAXdwBpeMitgBaRBVAIDmkP66+s5hIzn
C8LAm3j+T0Ueg/Js2GuiKrdJI66uh2bgrsEDBPXwv8mWJNEL6/7ZS6O0aUusIesM
NdfbH+hbPIb8Nzt9MejE/bwtdFv2EqiS63DLArJzxkXyRXEG6FUTIunc5QZvYXB5
KVw3Hskal8jGwtvsPEYcGQ/rUxzIXg0kol66iABnJD5Q5sJ+XOPNkR24JJ7Qp+U/
oM+IZE8YVza4leAji9BN6zJQhBjm19FQps+9vnVMr/gcz1qt9muAzJj8e4GsG0vO
eLVTna3irILm+SLVroQ4tEpPveGptINgsntxBzV8Gck/MlOaCBtFKnyKlsn7+Q1M
/kC9V4iWhTa1kkJxM6GTihP49Pf7vbr/bsMDLI34lIwGr0JWxUnKOsJdULtVZpyE
CLUIJ3kL9fTRzWtPChPxcsGgQjG36Usi9vrYFVJHshWco+730Lfn+7tAqdH5oN+a
pqVzrTbAryZskxE4ykNtYS630/RKokEIB1G4VDe6ByAzAaQh0fbKogNCoim1yg5M
ZvTm2DFKN29QObLLzphUKHxGig5lyOYXkx3Cx0Sa0Y3xfX06x63klvLB6j9wGHA5
A+HjlCem3Hu29zZom08NGZKPdhf0/Y2afImjmIxv+KbJF3ZGNhCVPnfiGCvd7I4B
eTgwNuRMwvWxBooJ5QJREAxRgRDlsK0x1lyYp+EtNdVrX4wTJNgPX69EH+FEfX8W
X1JSdAR0HeaSZxLQgAmkc7a0Ii7h2e9zeSQpKGo8gQEq6/Qd26DlTV9+DQcRWwZK
Th/s4CYxtymMutn8wGrLU12giJiOkZ4U3UezPxmiJjgxDIHh4buigIW1UA7QZGQE
Ac8GGmf+PnmdW19yWRRV/YlqE/NDoE3uIJrL9e6D6GzbCP9L1b2s1yiIJBHteLD5
KoZnIX5pUy+jUPU+ypzRWMd9ZTVSOVZMbsEhp1cyd1jhK2xh39y8famPzUJo4rPN
Hnq0Vbu+RpCHcQ5hOdV7p2obsGsjlKMSbyOk+X7UNKt7IeEIR8QxcKfQGZ6JrmyG
SvNoHL63gleyfmtY0SbXsgv6uXUbawWWlOMNYe6KUGoaXMyTUpxd/ejr9R64dqVv
hnQtWZSwSmkZLual4w+f27PdrruiZGERUOnyHcD+bnY2PaFMzV5MeJQFeyuc3/Oj
MdZfMaAMtGxOaH2d/+v4K20w08577sLLRO2MBR5uDW9GkihNZdhDrUSCE9GEHVz5
kCVbghkh1V9nHf+dmLXNnvmPSXQcHbpAtnYAaoT3H3nqCqWKCiUeLBKO/XmWVBvw
dci9oHZoFvwfxV7dkoZ9YK9q0rScoN11oEgvdrUHzONCNd9sBC5gKlsH9Wr0tEd4
Vo8WyjhAGZGivuvaydjkvVIoqiCzS0tGGpPPODGPiDkluIPjJCVYrOkWsHf+odS1
xoYmavS//CogINijfNrdhYvCraBSO4FNTEws35zfqN22+s4yHeZfgonezDXA6/nt
nAYr+bRb0poqMc5pHyBkdxh3GK+V6EIQUnbvYW/fRptPzLcM/+9VRClmxD4G4LVO
TsuL4DTiYYSHYTWov9iqmbB0/Zv/R+FWJBb2+4lbx7HOwx3SYZnWR2ZJ7OY8bSvf
xlVf30ylZY/IjbAez4A1oMHROaR9y4aMrlTuy0iqNE0hpUan/LtRBVLWzny9SVzJ
SmQyJ6Wn7rwklMy9vfqiuqAG9Ffb0mnPJ1vxX45GO3npy2BGjhRX/qvtQfJsEln3
IU4e7jF66vg75XZd9YGSWezCUFRYyog7RIN0HjUVg9Jq7Wz2cJDl70p9c1uS6kJN
2++ZOtzyUxFdXZkmBmaX9UMyeXmznfXWG/B4NhnEFzUI5NQwPg4eKupKQnp7kDVY
VC/mR4Qqe01Eo9Wn79I9U633DMR9fkGlvvLJLOMzxhHhQ0OBrYXGdk3CmRz17ktC
GTCIgw7r3oJtvN5vclYhj1L5XjaWZiyPUUxnax9rZyqKMc9rVyuNdUnv12+7JzWG
6tn+1GJgJiEA1diPBPxjCriD7qeGHBg/iCGWLZU1+OPlLjBlSsaWZ1GJrhDt/4Ai
8Wn2BMtfZXD9C2NyhDBbE95nADAdgLs4mDURuEmcL2/zNdl37Pmb4fcLWKv7Uwfr
6kNvVReHhc+aTlcgMTY8nHXlw0uXMZnfzWcyuMun/r+gMdXlhGqFVq0/p9Mlygx5
LXEq1B2kjmFwcqOcXIGtV7ArhF6jbTk1oeh2wOZJUyB60ctsLOI7Jqul+Me7M8dc
J6VTNAWYhXM97v+RNBYqGoFtB/V1n/7FhDJ4Hfn00qsDtiM2AtTw3JstUGx7737n
K9iuy5yEVPaQvramfg/rwNv2f91xfuVGt2RpqRZ43ZxQgcduGXxCy58DyKlVDB8i
X3cG7FcUBCKgloIExd8iNXs8GQeOvCVq+BmUi1K8YzT08MIUg0vTUWpHdxwxJGe2
ItVpsFcGjxGDh79BM2LscH32ANSXv9LJGOXMjUALhQgswE0ssx4rguSo7Dl+2X29
DDBYTufiKYMwIyIhzX3UARAgPaWu/Tgm39xA3CbJzYEmS9oezBQVvqAtq79M4g8U
O1PnD91AAyNmq3uRhTw8spEFayjtmQRQFWrnUZpnYq9jCZqvJwfjFGEehiYPDubu
ryMAZFfSpQOgYktPHkJT5YzGmymHmtavNDNKNbT2C5Iss3D343Te7upNGSHuMjd9
SwbAGuFgVl42g4kUy5D/Ed6/XXd0yByz6toyd4QBaw5yHps4ZARsHjyCEWctrrq2
9yHQpfeDfGyQ4Ps6kyzDcQ==
`pragma protect end_protected
