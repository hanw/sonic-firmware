��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z���+4eTc��:ώ�<^���_��I�ǡrP���o���(�O�ȋ�{꤉��a�I�SO��3��\��>�]�'U��2��Ս�eij2m���}�?�w Xa�PX�̈́��]M4�����.�v
���:
haa��n^�g�)��' L����N�˽��-�_���#��*���?�T�|����ز,�-�(g{R� ����2����'�ܠ��Ь"Fc�FZu�8J���A�YI�/�����*|�m�!�_��h�tã,N5nJ`�9FV��ػw��5O�Do��p6ET;��)��y�����пz�[���ԪQ�rB%���Q���X�����Ѐl��PHe	ǮJ�{Y���Ur)G��&F�Ř�ŋ���yq�V�Z�Ju;��By`}j7{�����q ��;p��x�K���8���6ĕ�Lߤ���';�B5|$8a�:�Wl~ �A|`^1��B�Kj:ټ *rV�%�qFQ̤�1���>�4�7��� �@*���E#����
_�-kʸ�o�Z"�����3q0{�lW!�͟h���w3)�⮬G�;.S���`*�j��ڝX��>{r�����-�%���7�"ܳ��傷���Z$U���ME"bW���.��Q,��J��G�9��Є��S?&�����,�@�@]�?��6VC��jb^����=v��V`]�Aq���:�S����Y�o��i�]�[Cס���PX�H*��a���Ed�na���ObB��1�[����HQoc=L�~�X`���e�D	Ղ�YC����WH=�-z}|��]br`�n;o3��R�[əO�@���3�O������[�ts	�;ĤR�Dj���dE��NN�U`gâ�2�3�����}�Ox����A�2C�G��j[���������P�/�p_�[oT���Z�#iT�l7��|�	s2ܸ"q�řl��>�>}^U�:JE���7�����j�r���ˇ�gh�pL9��((���Y��	��*��g�rHDAiWk<��WghC�{�p�4r�/���aj�d\e��BS�X�ka)~��B�u�BqC#r�F瘒��K1�L�2H��/~��g���Ln�qp��aV������kf[�@m�]��Y���x��M����2\dlNW?ַZG��d?0͇%�"ŋo�L��x�Q��J!G�e@�x�Ԍ��:��@\�Ny �k�X���%�k&i�kǻ��7XO8�ʁ��ATSC�쿖�1���s�ߌڿ�)�H���2=��_~M\�x�4�&�	���}���~��c���L��ǻ$����Ff�He�Хv�@��y�'�:�����>Fq��R�
H�7�}�`����]�]ؔK�>�a%Ǻ���0%���YLbdo���n�D@���:���}'�σ~�I�U�	������H�ؤ8-8����D0��4�}̶�.�a�W�yK�%�`�s�^'a����|N���w�$p�	�v�F�C }62C��R��	?CX�����x
�����$�jo�=Gs+W�H�����p�s(X�ρb�'K��^�m������Y,/����g9&A�M�`����M���:pf�4��L.���6u�m�͡ǃ���/K�,�����C�%��t& �o�6^rȸ,V�;>hr%��<��B��PT&�8��!,�x���'�nsKL��Y�~���j���	y"k�̩��:A�E�\�͋����(��kV���0u�z��"K.�?�H�N/�=2�_�V�%��ܔA-B���;s��/��
y�qޥ�tsj�a���r0W��qx���V"k&:>�oזU��a�F`	����$۲;C�Z_��a�0�^�j�\��Q �PhI�n�_M�ppm�򰓗A 	X�d�����_]�Y�a�*A
?MZH���Y6��'������j�����b6���"�2�{>�.�fY\��\��ߧ(Y������?;Ws�\8�ς�Ÿ�FT�!rSp�]]�"��5���R\1�J���C#���GS�0FX8wr�{ɰ~��+Ǉ+ ,;�@���|0��B7y0\��j�)�i|*�j�U�g(׎G�0O���9��W��ݠ���v�i)����5�������C ��US�-����k�A�p[ \�H��8i��a�����a��$/C�� ��fſ�?�C���WL�ݖi�B�Y��'*�G�R<�G�'�h�;�����@
B��d�p������ڃ�YT")��]khS�Mp�w���G �7)�j��7)	+ ��:�D��+�^/�KKH�$2jyx�����pL�ox?$yCkn�ƻ;@�.+��u�t����e՛�6/b��>�2�o" ��	ҏ,g�幟UPE�끔�呸�쉭4
=��)�Z��!����߳�#[4��}V?�U�؀��C0-P餦0�lΡ��Wl���݁�R�1�c�-՟�W.�}��.�1 � '��