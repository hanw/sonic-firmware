��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���/���K}W��v�!��~V �qc�H_\�O<�a�S�*qI�4�gp|���ɞ��}b�
���~�񕵑S��o��v�6�Z��2��z��O'-���
�!L�������a���C��4l���H��:��ŉڰ�ZΟ�u�"�\���/�{a�p����l����=.Ndd�/���x���M�~��N��f[k��a6�;�q�Ep�J �N���B����?CC5��>ϵbV\���}F��ݗ�զ8U�0��hV���3S�!��yl��e���4>����bv��_[fb�i��Nh�}̞]8���@z�7��Z�I�;y�x�A��pɋ"!�x���I�7�*&BթJ�O�z��p&�q����֘TfY��Cq͙s��J#����D޲M��Pd1��Ng2�x2u�����F������%#B��y����R��3�xM�K��>��?��v8'*���d����p�]���{h,��p��H�x�� R��t�O������n�`vo:e-僀zCy���,��=1��ʨ#���~j`�+��Qņ���Ҵ%��IF��XWR����Y*�l��C���'���L+uɵ���s��O���SB���]�4@`!0*����ˑ� ����$q�o�1�<�}��C��nmi�k�N3	�X�*����D݇�q z��$�.������K�g�����8��h�I�1�b7��1�+�'���{:_#
���ɠ8������sf�`;#X��� إ�s:ŸRu���~�H��S��9�HGC1�U㞐.S��&q��#�p��P`-5[��G��ƞ�Sfl ؍48�����v���`|-e�A�x�w]��e#�WO5��'�Λ.@R��P�l؏��ɢ0'N����%�7I"�V�W�d��L�²
;.Qj��F1�|�
֙���͜�Éǰ^��2P��N����4Y�k�����B����5��FBv���J�A�9��x�U贉�C�x��W�&�k�c�fY#�QzʏJ��c�(s�ë♒�(���C<�Ψ���'m��&bb�W휔������'rvMe3,0O{,��]��hu�4@�Y�]�����0���H�vx�_�jf�*Ѧ-�f]�M�����xdv=�X�|������JS�>�KM��]�T�C+c�o<�F(�7"^+�	 ��b�<�H�tg�?0E1����q���9�9�Q2���X}�y�k��+P��x;aP��QkL+�Z�U��	+@�@���
�
$
>����˵�>#9�u���up�#�����v<q�і.E�w��zu:��)����r��-tɈ_ � �Gi��8�'���������(P�?7Ê��d��Ū��~lDn5���e��wTb�/���.���{�4�P�� "C	�������?�l��¨�uW���Gl��\pQd��m�ϊ"ndlbɡ����6�*��\U�ɵ����_$,���g��
RA�l�x�x"�F*(x.:�B�,�l��:�(��p5䷱�o-_�i2�[:�aD�� �{q�;��'�i|�P�@f:��z�*^B�;�J"a}�T_X03��`r.r��0���`3�4I�Z/�iK���=qk�nG[�u��SCO<�2��,g"i8��90���g��#+s_%
Z���o��3cŸ{�Jo�}�.��cv	̇��	O$U���'pis�PV���B�Qr\�� ���� [�ȱ㌢��x4�4�-�z���M"�*�j�v�0S�³n������	9��0n �p ��r����|�����w0مI�����Sy3����=��:>䷡�C��'�p�KP��� ��P���/�2q��)����J�;X�iX�j#gݙ��Xl�e���zp����J:���	 ���!|���z�O3<�f�fO���_�^㺸�Ո;�%�)�p^~y�2�%_�]��$�x�=�5�]��_P`�H3Vr"A9��^2�w|��7��0K�U}�2� �]eFm|�sY��}��"a #=)�O���!G�j�r"�>^������'�e�WǪ ���Pӯo@^9���m��rFS�j�P�p��:��� �����:�?�8�i���W��"	���a�u��q�37��������#�Z�Q�d����tS	 M����6c�Es��T�xJ�)�7 du�gMmSm�Q���ZZJ�a��9��9�6.�Ir��ag�d�i��N��BN���h�#̛���X��V�<F����ّ�0�w��Dx^x����[F�.��;:���Z�[s�ᇭSo�[�+V�3�U���/�?�c2)���9�'*�F��wP�:0$�Ȟ��˾���J>�&K�k��W5k���y��lE����v��1z��� $�Z�e{�� ����)��΍Bi�sIi��(T�_S�'u��Mx�(�����\���P�;:�L�4����!Kv��T������#����l��Ro���,�n����o�r9�	�'|�(ȭ�9�06'�{������+�	�Ǐ\�#��ԓ�=��eS���� 4�&�����C�s�qHd�"�!��\Y�4F_ <�AY�����H���B��-�¿�TA�NU�*p!�!��	S
��Ƙb�	���f���
P��*�M���G�+��	U|3��n��i��*>/"���-gup���+�S�)Χ��6����:�3��N Yu!�0���ݩ��K��2+HgcS�����l����p��XJ���!�F�&\M��a��.r���z�IՈ�hK ��Y!���?�dɒ�l*e2P��)͎��uP�u=���b]+&Z��ɻ�,�+��>  ����lcrG�]8i,I����vy�sC\��AN|�GgGkE#@��*���7��H��;�>U/?�`��,&������7"̍�4�ے�<��r�(\{�I8EEۺfz������i�w��������=�h��ͱ��^	%J[^]q�WB�dt��-�+*��HGA��g�HwJm�˛�AJ�3y�3\=��T)wȩR\����˯k������"8��2R2�Hn��j�6P��)o��l� 琟"|^��2��LSJ�zkF�y�.�(j�Ms@(EFU����,�'��H�Tb�DvL��E�F6w��h[�祅&Ϣ.��kGu�������U�!�hEi�>70|ߤp`�62�3�����j<���8���^ڸ���Ǵ�B:�o&��c4�jm揊j:b����S>���B�-�3~}���^@��5L^��x Ҝ8�y@!�g���z���B�&g�S�Jn�*<�V!�yz�^A��Mq��/���O�M~��ndC�8��zu�3Y�?������w�^;1�8�4_^���H��G	��Cv[�����^W����.f������͘=�f�#�YS"'��T��8D;izR�)��:m�a���� c�H�&��v ɇ�0>��W�q��>�v������"�,���U�,��>��h���R@��ǡ6.�S��f�G�"-� �1�N��dڻ����%ְ�}�w�m8*]�E�[� �T=&r�8�h����;�J���y��b��zd���ԵȋF�ay���Z1G&�pI{��3���?�U^u6�au���X�Z6̓��?(� ׹�����ěl�0A���q�����>Z<ҹ
�صThI�un�7��8�����|�YF5�ʼ�D�*&p}XF֝}�NF�����X6���s�NBAp�=��
�4x��'��7of���W[\Rn���bt��* �_0�Z)�:>˔ ��P�c�?��c��0`��D"'a�2��3������]�D?3.�$�T���>e��v�$n�Z�kԙ���&2�/��-�~sG�(	��N/&��ku�EF�>��Gtc�$[�Y ��Lj�0Y�����'6#��#�q��
�/���B�D����K���vw��/��؏Y�h+��R���f����`Ŧ`�&�Y$�g���pD:�ۯW�}�J��{�<�r�J���@("�+,ҏ��/Wd}}Q��42b�<�h��6�}ޣ�8�WTi��S�^�K̒ƅ���ß������ �����+�d��T�ϲ��[�f[�����6�&�z.0���Yl��8O����cAE8;t��r���k'�.�#&��q+��������Ǉ�fnй<�
�G�H����6�#m)�^�����3&+�H���5�# t3/w_� XY�i�hb��me[��hq���a�i�`iRH�5�?6����i?�$_0,hzq��� �v��+y���y�<.�u�B���-��|{��n�A��?<�S�����Rܖ�u����Cɻ։4��y1Vީ.č�E��*aa����)}����t�D��&Ǻe'(�HW��;W�>T��[����l�
��p��A�?{ȅE��dF=������+Q�r�����Hi�4n8��+y�^k��ua���;|��3(�Ž����Y���u[K=젲Uթ���V|�1�8Ua���G���]g���s�`��TL�"j���O�b)�>dF���h��<�ߤf���j�����������VBw�ҸS��\�IT\���|���&]A2�b�.D��5���88�H�.��4TWK���1>s�}�@�ƨ�����D~�|�u�ձ8�ū\�C	a��̤ge;N�*���y*�z��Y��T����5�Ld��Hl���=��,�U�1��rl����&.PJ��Ǭ�,�7*����bt�I�V�#�,���S�"�c�gN_��ʗ&������^�&��)�(����w[�َ.��K���\AX�u8�vt��2������b��@\F~5Or$Z �	��i�E74��~�T���m�;)c��)s��ڜ��Op����"������U�R���qv_����?k��Z獒��o��G�Ȧ"��I�)�Ft_�M����|�rf��J�Ps������+�,6�� ���gιKGk��D�b�N�`��"nᎭu/tV�-_65,))9����#@ _v�̘~��\�?O�|I��!B��z����)5�����F�bX�r�?���<���
SZk'f8�)C]ZP\�p!9^"�a孂�9��S6�l(�É�kJy�夽���o�ќ�@��:T�C8ͮ�Z�E�3;3�Yb�)3}�P^+m�G�>��=�r1�k�}����j���x�`!~���`��މ�e+��F��^�Bѡ��(����Wy���G�k�=���҆����q�S=a�nIjW�3�k�`�wV|_F��.9f�E�	d�ȆpB�~4�N{%�TT!Ip�^*`�h���K�+���,Km���f �B���S�Y;�	�Bw�S�`,ل-�	��y������W�x��f��:������<�A������hϱnf���=t�ґ�R��3���M^*m��$�[�cZ��l*�e?\�Af�=f*����z��^�4��9�����zQ� }
����oP�l��n�Ϡh5u�|t�	�e���ծF�b�y��9�Y�]�=T��Z�wj���w��ɐ�m���Kh���+)PC�X*�&GQY2n�@G�:�LejY��3'�\��YU�48�Y{���D5'�5��BƮKP��uV�q���>T)��>-���$-���9V�f���%h�-���'��2����g$�wi||R:Rm��
����|\�6#R��/Oyn��p帚ȣ5���R?E"���d\�/�օ���c��r�g��V�إG��|1��6m�V�l�NOwD<ڄ��;	��hL�d"���X�6�I�w�姜�t�i�j�{؀�[B�������-�1�K��Ws��đ�5��TAE�<���LZ�ˡ� ��ߛ��]�\�K��a�'_�rM�̊Ǘţ���˟�����E�����Vr�qXnU��Vƀ�ob�R3�車wXq���\G	���\ �L/�ֿ�m��-	^%�١t������>�F=R�R�����B�SR
�S����?���Z��t����?�`�V�����խ�� @.H�T���<G\6��`M�6��� }�K�r�ժF�>i]Y��75�;֛aҳ�>��{e��57rX���x0F��$�#��n~�	���C��-��~�-�(âGcZ߂���o/���:��S����M��VI���y���_�{��ښ�4cr�P�Q(��s��UJ�M�e>edoe���&h���nP{LN�D�pZp�M�B]��f�u��g�Q����/kL�fh������4����	�|����4s��PfF|�.M����
9����_D[=�d���p)�3�tW}J�c%��w��)�ʞ��Cn�Y�Q��+�R�1��9��� �ُ�t0�f�q��F �C�Lh�?���bb�ʥ���W���7�I�)�A|{e"�����`ͮ;����B)+B\�ڽs<��o~v�r��w{~���S^�U˾��|�%�N�Ub�V8d�:M��N�TV~yFh� �4���GT�+����~��mɊ�~[%����Ki$���6�Ec�7<�rf�7.S��9��A����?Ju�^�56&��,�+���x6��GtG/+��|A�)"���j��U�I�׾|]b�E欟���{LàB>�{�����ґ�'�c�i4�,�N&���"���|+{B�*g��q�P��U�'zڧ�5�.�=�4���6�dXw�����8r���芧�z,�+�pb���Q�h�	�sJ�n}K���J�*�dg��sUJ��*�kG�~7ۿ�F~s�$�6'=oAʙ�K�a���e�&��"{@;�Pn8�����M`}[��Obt`L��￑|������i0�O�A��I�����=�(R�A��������}�ia"I���17�o5��3�5�ޥh���f���N�^�T�� ���y�J��c��ba�[4�!��2���M�����
rn��V])M�N��5���`4;Փ!*5���!-��phD-go��]���w�D >5	��99K�!�.�l|��9j�g7�FRl���9�C/� 6��5D
��*L������B� �v�Q@�n�����&����;��o0�s�9v:	�ԣ�j��������.<�$큞p��ܵ��F#�`\#k��ʁ$�l|>�b�d���ځ��[b�,ҿP�b{�2qp����j���Yd$��?@V�?��xw�l+����mTAD�Nٛ�k.f�f�B���#�YC���`x_���{��_[��~u}ϲ��v�{��U�b��dz|�w�n��Q���ܡ�5��&QM�ΰ+������؍y�N��M*�d��Am�y��8F+s�����'e6[k�l�^�o�c^��rg�MyH� ��B"�OR�B�Ӛ�,��j�w�Ш�eWb�%G[��p5������i��M���t�w��J�} �z~/����ۦ,�ʹH��k�	�'��q��?
rF���Ǥ�R���p���ڼ��_k(��<uafjp�.���<U����6JB�c��8/�S�֪���:��5����.��T�������Y[�l\�}^3}8�W�XDt�M3}���m	
�=���YB���y���QYet���O�ɟ-�(&`%�(��_�T�"����I�4R��(?{�sx����A ĞM�_���S�[�M�LZH���B:�򩢾ֳ8-��u��B�SZ�3���7��1�t�rղ��"g�8�~:,D�wʽ�-�eu��_��Wø�րs�T�A���i��_ȨO#ǵ���v��