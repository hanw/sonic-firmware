// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
paJbLnYkDthcAwxQVC49OLHXo7K9Uh0UVrF9BNacGFnnyjY6md2Q7FXMhjBnbfhV
z1Pnln+vpd5RybQZoaw+2OBRRXJ2QXa4ZHxhFvVdMKHj0mcpFVklafQOxBc4grv7
DkVkdBHI78gz/RhpN4AoKXGIx4EgKPIvqdfoTwbXXA0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3424)
4siB+3GtvMMAwZGTKdnJBd70oU/7fpv/qVX5aCg0gT0gGAuTVP+ffsvhQAMLZ96E
YozNwHa04czWCwUI/6en2sbe2vW5rehExaYkZ5MCa4zQUiJjCUqG9uLVr/bI+3HO
D24G/3m3vgAFlTv6w2zeX+DBi7hN7H1OvtDi+U8EziSMMIsGIUbLhb+jcVMX1mW2
RsIOqXFEz5I4eHdnaOpu3z8LqCFNDrbbvfEfheViSeIWhQFt2yUtJRyBVb/duJHv
BXc02jlVWLAPWZPEnJBN+qPUHDMDxpnhnF2Q9UTE+xXRUa3GATEmz3k6RnLdLGBC
HrdnIuIN8h++/HDWD4pUucMEwWW1WbmQFVrk37BALcWn9eb21dxZjlrjCIP686Wf
+FGnMNYp78f+M1YFOXugpiGq3TWJvBDRpUCl0T8VyzxIgWE1O6etTkGwgy5uSzXy
V2VxvasVqca49bjIxN4wYJS1b9zWPGcrpZn4CX9vMMhJJMfZMnD0ABOTghiMmYoP
x3fpRhYe5hemiMQzWWhUY4xN8NyKshTlJdsD9Dqb6A2wg2V5d8N+e4MvZwJ2S7WP
v6w7nhPcS9B2pKnCeMQxHnWBBrSt6Tt8WtSaJZ6L2SoBY1NbRYj6iG0eQjictpAb
CBZsKetbgzn8zBdeSEs3ZJRdka7BCKv1ya62/o/73omF69Dl9fdwrXst4UwO9J1G
gpvgK3qkewXlIkrtOsua2LPTvNcclfaAIbTGrXa8G6qU0Q8WjwWOekyty9smctMs
j5yjA95mT0UliRRGAzIodcFW4lE+7f69duYepyZqfw4WuCOcnthOdVwSSjn6bDRc
k3DytlC3wviBQGtWpfLRBhWV9ru/Yju+ZjVLBGAlJwolI6V2clZKExY+1Pdudqki
CZAdrMJTuK5THpWk3nc+4c6zlPTEXazjU/95tYDaPSRTvAQRisTDLGR7r9Lhv789
6EbE6g8WEO/vSImKIWErWa/sANylkO8HsPtavSF9s1G2eRjRNkU9RkK6dRyLyhQg
4+OZU338Lhjjr62BjKq3cOteBMXJXShVJoDqhGNDN5JxXRkH5KddNxaxRvkCErIk
CQghjrateyVT4j8GYA3Y7wV+JuycjstDpbo+7ayL1t55lh/amTfI4X/JlyHuIK4n
OfgzMGhteJEVlKU+SzJNWmARNbemGX49/bq6lZo4k3OaNcW2IO9JNhEHuKkwfPMu
wI0rxmGzg5eK4gwznl0NfuO+S8mZ2sKWSGE/gXOUPpepZUZctAvXbt0uo7QnvEgm
VqSh5eNn/Mhq7rtzJjZOOebb6zsM/3Pa538TPn1X5LnLL4ywdXiWIkpnkqsB/XJt
olhP53wPX27HddPNYeDpHI5WvJXsslUT1I3V11/yo3L+bPuyL27k0xNohfbQFoZ9
/Wa+sMdZ5UYO7zYmSihtb7v6E3dXg9/zfrazD1yXAb0JwGdpxWn31STVje7NQLdS
01DjoLeo/hybfa3Mi12XHxpIKWaE/1AriQWt7W7b1lipSHMwKi/sFRpBbJfu1vIU
E9j99z6vnYEBZgbt5IjPOUyvHfFHBNVWbQq1RjPn6P8VJDWcRFfb39v3J+g7SK5e
1WgnNDt9UJW3urqFMbqvz0F9Lr+rkVYqpPkK0JKLGwv9FFq5Ohidkh8trfaylkPO
Rt8UqQqlfhv6gzY6hGm8VcTUYStOh3GkEqotEIBA43g+q53VKmb1VHSOwQqE3q6O
8KikIJOv+3nJydZWs0p0iN9OkfSpRFQOkcMYQ798V96hY4NMUmx1PRAtQ3zLErxE
gGrq8+vryIB1S0zkUpMH96EIhEd+4i93Q6wpcYFPEec8b9m/DEtH/J1fYrbNEmWi
uRtc5ykNWR+/NnNzRfUxUsKtpMLqI/1tF32Dc2yC50I83DpYL/hEZd+P+F2E+s9s
ZP0xOFKpd/avZUusuVMcb9omsWevbItThOCMDskK39VAM8kVqZ1avSKQdK4Sbwk8
MWYlV2MTAwTQQNHyyQJVckwPNrolVag3TM9s+AyBFeltRMIuz4zB7dZ0QPJN5hL1
iFaXFag3Pbgp7DriKN2LxpD1jb+oNRHiT8wK6Ysg5QWPNvGfZP90iFmXgX8NOR6R
JO0GTjyXqi6VlpC2D72+j7AUQFb/Q2Y9tYeXeyTEhHlbKWaNn1spNw14upLMAB4F
y1cO7ygDRaYXhbRBL9ZduQ1QuiRNUdguEiYlW8BXaUWh4pXq4Ryp0N1zKPSee1Eq
G3ynMHOtlenOMGuj/uXKHHX7soUW6yNMoOCUGCM5zwPR9RaqZpkxgmpaaLiYH5Es
RjAbAX83VE2rLEMenTa3DwZDKNI9ZrFWIv+/83IXu/IQyktB+FCubfKbM0vZjMi9
oePxjTzj1oZvLxl4+1SsMyeoEh/fuFd/vzCK5WBm1Ml9T+NTacub4vzD21ccX4VE
IApJWFbNmc1JnO1pKDeku0t1M+VJ8VbYi+H9kb6ceRdS44uA5/pPdCyDXjJA1lyj
3fGI5pBzr0JhhxcbE9j9Ac7hDrTFmufvbd5fLiKmvpJ0uY9lRRRVzN+sLYAB8JdX
mMv7FG1QVX7VDd3m9+Om6vcrUg6QxgLmIMpNdBjc5BrRiigr3/GnoQrGdyshtFCe
XfmydHTgzPBAz1ET5rHD+DV6mlXqpVcTmCvG2NWLyupBYGnhbiTGcC/x+MtnbVQa
rYiGjPSsWZL+t8yt4y7CBN/4C5Jfc0w0r7FQyF5qSN0m6kXH99jCCCaDOtJn966r
wGluR/LKO0wBZauT26XbTC3vzeIZG3u4KJmC3zsWOX4ZNjW4UnInue/lapmTieWP
g+mZEWqqeQjge9sikqkI5RgZhS/WxiHDwm2imi0rKd9hOaZl6mpk3NKxeSPloWvA
LqJMuWKBPaNw56JVcjFuBIgWNigH4MmcjF2XS2hdxCsYeKqoOYQhtqIw9FV/jpwM
d41iQVgb/WrjglCkLaq32pkmuYaoTlLr32aNE4UOMNNAeElW+qniuq+VRCku7iq5
irmiK7kxrt+HZT2sxvYybRAKjFG5OFe7Yq+3q3SeMqMJ4pu6AuAvL8eKFoudeWFX
IFbw1PRfFBblo7aY0xthFqcrjCetEB+qVvZEaqyRf5Wq65swLe2Pmq4p7tH0wXEH
ljyb9fvThnf7+acjQCGWY9FA67Bl1BHtiPkpwPFt4T8nLvHXNHXf67JkoN/H4fLk
KBxHcvfZZeYw2980p3B+wUEfTOQrDIuWDNqup8Xy2hvh1ovL4WZcG0f6JE/2BGs8
bF1z8xbGnioHCzoawOmidn3qwErOokxMtY2itDKEP+ky6nye1zyhXz42Zt6cn1ow
nFMD1il7QZqiogttZJIRl3aCMazSiyx3CEObb1DH9POMWXkV27TvumAEIKhgZBbN
FImsuNerBa+9U1js1JfE1PKTwSFQhRShjWbNzJKAzeANTXhj/ZyI0pZB+AEb+DYH
HCoNdOxESLDjSYlFrFvGtG15UdnTo9Pz+wWmNi1eaZ8IQBOZsCPIDnLeW+a/ZCdJ
Y1nWKw7LXg8tz7me8kKgGWwhnoAL+uRgTYD3hPjmwXtJM/Vo8T9cw8PO3w9uPLLw
P9REhmtfbYMQqS0Ovy/22h+5ruzgtfxv33PKsDNMJSBgplAVGv7zkArObLI1EtYZ
2T5UgDIC0n3ZKHAj0zcV6SHBT2DnLMNwEA5D7FGAnwavwsHrIqZMyqH5PDndw1EJ
cRxqilqS2bkpjlJSbac6o+eFCQASOBqDfhpryqjiFaAILiYtIeVoRx18EmqASbdT
J8jkBn/mCL15u27VyO/8K6xaCE4a6RpNkslbs5R5jBE3suPA3Edk7ryc/tq7sOJL
8u64sqO00D+q8rl6aHSn4Od3Z9XBgM6fEuX826aDToKQJz4JKThLGDfpdksYSNSG
resNvnFQc9YC3oDHcVgSgFHt9azJ5WbHWyvAAO6fJULRSHHFYwiTzaAJy6e32hfy
gEZ32/wRHMSaC3+XqwO/6TaqmmodRlYiYHs8zOq5FNTp9Kni3zNZRNwesfxaPP9g
M+30MZRYYfABNWxi8/X71/pnHo6C2BQQiU9Qj6Z7K3d6xF+/zoHvP6kIAQzVcQbE
+UChXVULrKz5BFTZnw7adbuoAdL/dBpvTVsaldvXzPco8h918r9Idtk1WLbHEOkw
Hy1PzmDY+NJLa9c7I51Yjxleco41l3NPlPoGiSX5CDiUvXMk4f/GbL7zR0rDxfaw
Aubh+bIEQyUjuE3fTbjcPalzvexiUGHuj9ZVAXbtIe3xuueFtB7MGSQgKtE1iCgB
CI0I9T+TLR+SvHB5GJ1AYU9pxx90Mg/VLHI1lGH9Per8YeWQIcpyE3G3u1ZXV64d
f4+zfuV6B5GT7BQu2JTTMbRmeyxoJLLQnz5QE9p/GbD1kSGXxy3wpWsKB9qBkRd7
viu88k+jd41odsw9IO/KBZAtkHRRhX6gsM6Tcv1VUWXtDHHoX50TRURoVhvzjZeP
ectfKlxsGRXgODcGYGkIUqlkCNtI9WNr33nzdbscrV+rhSGazo6emvQNExZv1/yd
nLvEGopKb+v7eIt+EFy0KA==
`pragma protect end_protected
