��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z�_������L��|���ι\Y4Q�f�B,�A��\� ��鳍I����vTk��n�31ЉG�Em����.�x�v�����C�A�n�eH� (�g���ܒ�O@�s����Օ]�$��*�U������[�7Cc����#4��:�����N��l'
�\��t�t��j1��O�o�9Ulo�������F�����{�J2�>��Ϟ��s�E�d������ZN��'e�͢i�J�`7��mEY���[6�]WQ��BՈ�M�Ց��-���anf�рE�$Bg�ҚrF\�:`w�Z]F�ar��,��eю��ז���ε�ۻ��1L�q��i[J���lԷe2�L�M����C�t �4l8��'*3Z��$�9]]�X�V��,���i���Eq��jKc��t �f�T�8��}؂�C��S���S�[M�6�*��(V����uA�𿁎���xo>& �-H>m�*��@:O!"��N�Ǡ��m\�����9 BɈF5NKى��1MDGԞ��L�^�%���桉�Ql�������0uXyd��i������ �29,Z9��j��ݲ�V�OL�J��B���B�{���������_�&.ص�>V��5��h$�@qqމ<�r�/���H���8SZ��M��2Z;|4,/�����Nn�?��07�l(O�
�|'B�3������'Xhd%Kkt�������jqz�窖񦿢�ԘJ\�.�5/@*�2Qo8�w�%�������~;)�,Kz�bns�HM���̠�7�/92�����g�u�=���K#:j�בX����`���%������9&��%"�,��hd�9Z�s_['4omK�������Sh�i���ܒI�;7mԔ$y�:�M�󁰒��H��g4�p=�2G�3�4��Q����ej�]B���ty�x��9��/[H�4KH�:[q�aC�5\l�ه���-�J�y��q�z�����bL`F{f���FYw�tپn��=�ν�To�ٚd7�g��'�C����Xd�
Alk�Vg=X{�����~���uJ�+/���U:��4$$��N�ɉgm��T�|h���b�W��p��ȳ`]�m� 6��I�����=-�k�����D�mx�{����3�Y�:t泐�;{���75��Q"��u��=j.D;	$9z�L�O%��~cFV�#P��t�}{� 9�#��S�����A��[�g�hdP��{��g����!��~���Q��o��nʎd/h6��B��`�����w�4��e�� ��o�-Y8���f�)�j�dץ��'�@�rx�0"��	��8訿4Ϥ)'��[�{ۡXK�H�)���1����Y���z��B{�#�i_gz,}"�2��˷�Ʋر{�v�	�1Yɂ8s:�?j)�ݮx��L|Վ^(�c���*��MJ��7��j<jp�_D0e_E�Fxp(��BXt�e�e��\4��ځs�<�c��3��3��'��9	��	��uUz�c�Z�4�JX����b�G뎫�Gd!��t�����[�V��9+|����%>
��������)�W\���N����r�k��p��){��υ_�2���d�����*4�p�-���A��Č4w���	�4����3���|(D�p��B�$t�xD-��T<� mk������]`�-��8Ko�;{���β�k��9�����\�޴����=S<�Ԩ�Tu£D������⠓�BL�껵ʋ��4by?}:&�٬��+U���p��U�墶�!秭)�/�f���mN�& �����&ܩ�:��L�t��j-֓��#���9�ƀ|�5^��|���pb}����W��@2���bG�U_�@��S��:z�BP�A/~��	m�?����[GV�VU��=�Y�ׂ���^A��S���<��I��]�^��CB�����ǖ��_MH�l���N0Ā�+��#��)?|��V�a)�V#�<��~�bO���$��M;��2N�clUM:�!�����cq�3�r��]����驮ld4����},(��6^�Hv!�h�yi*;��AHd�,{�#��_�e��
X<����K�h[$�th����U�R�P(K�bF-��na/V3v�$)-���`���u��,Bg�}���O��ԘU�U�{E�A���!،��ݚ����N1ƴ�jlF������3�� �~��y-��k|7��)�S�g�j�N��Z��"��}��X���4}�+�v�F�/��'\=��+���>�g����>�����Sڬ��������P�����JM�s9^�T���.�w�d���y#��zƓ�!��?�jK�=<n<���
Q�;���(5Xa���=�������J��]me]�8I�"CMt<<�<yY{��R�>���ѳ�W�9'��L�\�n�|
wQ��$��4P i4�]р���	�� �9g\z��N4��L
J��8�H�ej$w��3'{�����L�i	�[(�y���A�.Y#LƋG`�]���X���X�� ��1���J=J-��Wek�	ư�ю�`�!Nu`��L,��P�n	N�qz�U���`�8ĭ�b�;�N�lx)6�*��Ј����?�u��o�槄�^��錉+Λ�Cμ	?~��DI�mq�����xr��}�U�w����Si�mYU��A�A� ���Y��q���뜽N�>�d0��Zk7�$?����K�`���������jՉ��U���j9	�3!y�-\U�PZF���w4^�E�i���Y6�=���j����B��V��\i ��Rr`�%��b#��x�^�D;�*�<W�]�i��R��GI��[�"��7�z�6�9ڻu&/]4'J��'x�2=0z]Z�F���(G�jEP�y��H�Y��f�9�e�l�l�_r�	����ɉ��P󩞪�&�3hC�P��1��hr��2��(�T����W�P¹�^�HAu=�$��ie���?�<c��br�g�f;���,�����f�N9^��(�C4��Q��9`o"�l���.��]+Z����GS�r�d�E^�p�>�' �g+dͦQ�1�5>��X�~�����ZX�If+3�QN����ma�����xpdR=즏�D>/L7��𣺍������D��c3~���3�i����/�O�pY�;�����[�V�M�fш̻�?
m�}3��e����@��������CS��4�j1�!��h�{3,꓂%\�n@� �~C#Ӫ���Jk���j��#c�n6'�1�����-9�Y���7l�#��@�����T�e8?p�R��k����`���s���u���BJfY�:IOd�%&r�ޢ!\um�6u(��Y���ՔX�d���g
�V���9�{`8P7����v�,)����+�a&���J�(�hr�Q���R�l���0�/���1>���&=�J�UgDR��F!����v��a����A�8n��J�\��.�([O�"�'�j`��M��)U������9lͻ3[�[≂|l���@�!�l�
�E,�X��TFˑR'\[�{��J��u
@g�//H��6;�o� �s����ŵ[�+ʯ`0���:݀�&Q�_�ȕu���{�Z��yGWL���?���W�	`�a�ma�_��-+�(�\���$��A9����l��|�3�M�` ��k�{F��8c���W�G\v�5/�y�)a�'Il����bUZ���W��@��Q�^4K�8c��i]J.�;�j\p�+��Hu�)��?���F���V(�XlB_͝����)��">��_��#R��v��}�Q=J"'c�`�*=��H�'!g*� 78�q��.�~�*�ٻ0���(���H�g�Kh������b@��)� c""\�w������Ǹ kG���Y Gq���Q��pv��5�hP
A<VG��)X\���	"wr��ɦ:�@o7Z�)�!�i�#W���dv;4���1��'��x�(����R%%�������yF��D��A�CmƦE�����8E�m�e5��6n�W�����۰ytG����<`��b{�O%j�,(u�w��6�6EП��o���24�\P� rn����h�:j(�:m�w�!���a�|�DX��E-'�a�v!qX�"j*��4�Z�3O^d�e�r��[G�NLe�z'�_�7ml{8惻���(Rč�r\|q�F� �qS3#N�8�q���S�Fj2���{K���\�BAὧ�	l�f+�M���f A���xu�"��!D�*�q�آ �W�b]r�7�d�;�8��m�{�8�+��kT��5|��(�>��e�	��k`�!'��o�+&xG�ni˂�|�6�Ε�|;�S���T�:"�á���ᶭ��ٱ1qTU���"��S��cg[F�w_��:��8.��)ƽ�AR�!����H]3�L�c�r���]ṙ�P|^՟p��xޖF�N�j��E�!'-LQ���+q�nI2
T��g?vo"�պ~6B?�FQB��˖������aT	�,���^l	���[��x=�rdE�s��^2�7SA2�T�����*":ч�޻:D��FG� @�#s�k�+Q^*�߀�^�Q�%���}��F�$����A�V��c�{N��,���	����d#4o��EԦU%g��xK���0.�iX`K_���|_�F���6����l�SwV9ZUr���Qݱ,�~ı&�wE}�nK��(�4Z;v�@� �$RQW�|+���t��W��í��
[���@���ͺ��X��<��2��J����X�p��- p񸅢@D�\E*`�����<���[YR�R
�^�2��i���!�]B�hasU }�\��g��"G.YhjE �ca$�[H�;����j!��hd��<5OZ����$�om4,k�Ec��,-� o���iH��V�[~,Ԯ>�r�y���|�S�:D A���
��+�>Q,tI|�����;l���Y��\�5�mLa(�����NS&DE!�x�ߗ׹А�2oyW}p�8)�מ�[��6v,�	��7,��Ɲ8!�X����`}�N�9�ǮY��z��Zl+�3&%�lt��s��V	�:��>�+bҚq��,�72	Q��;�t��?��&����̈�Y�O(bB�VG�Ԛ��G^вe,��Q�IP��sG;u��F;#�V�A�@�����z	�W7 ������*&<vȻ߁�e�~�$�H�5l0R��>_?�����,f��U2��3f��u�;&�
X?�L�c-;G�۫�{j��n]���Ԃc>����X$��2j?�Q���a�\=�����:�xLgmu�^q��j�b:�xy�6G���A�'�oշ0��Vz� 
��SX.��=�;c�t���m��똅B�3x�<�T,��3؋�7ͯ�g���'����|����H�S���z���oEJ+�Fq<XD����$ȼn��~|+�G l��*I܊��G���?���T$G�ٌ��x'Y�\&���.}��͉�jہ��C���ԙ�=�nu�wڟ�S9�D뻒���z%�����?�����p��fg�����2�eDs�K�6v:aw9�dhm�O�b9�:��U�y$4� ^��e�`�5�pH��g����- XT���6���vqX2��@�՞q1c��	���.�g >���_�N�GH�Awg�|�m��J�7(����Sz��) L
��"xB�S6����؍�8Y���fa�b�gNk5vvLF(�0�y�ʌ��S��*��E�eC0����>qT����L��Ý�_~���9�U�KiG��g����m�B9}�[N┺a~?��]��3~���T����glj�H����&�f�O�����.]�9���:�Uc�;�������_��gU�b^�_����J���c2c���&l(h�������Ev� ���Q��9/�3��g�ú><�HyRq׬}���yϪG�y�r2�ʲcu�K�;p)@�����yZ����m7r�dr��0��Jj��h�T�=��n|h�#Dv�����f�J����jc�Ƨ�����~��5n����;�,���qkQ )���:�p�A�}q�xA�����\-hKP�<��&��AGh�;r�Ak����s�c�骷��ȱP��`APY`�~��H��L���~N-����T6��P)]tXo����Q������9�q�G���@���@dc��Q�gdZ�~��=�=���m�;7�8�g���=V��It�@[�@>�$�Rz��בUyd�������J�|x
�2��C��{�\[����q������n���HL���:�(�3�<F�-�����qa�����lao$�����)�������ӅH<䒰�e�=!z3����I:@?�Ȓ���/�8��=j؞��Jmv�>P����	�n0/o�0$7iO�Q��� ��D1I9�_\�tB�6�g������A2���X�|��Ym]9h��X&%K����*��w�˧�mҺ_8����� >R`� ��5�;g�
�����b^�&�HA�|��NLa�Y��z���2�?�cӦ�p"RQwWd��q���M���a���ES�yh��ӫPruh��ckp��a�kw}57���j���^DPT���G�6P(��,�&�~q�x�؃�NN��N�����wuK�k���w<Ǫ{A��zox�!/q	�A�k'S�h������䬖6��mܼ�Q���s�P_�};�P���-@��[\ ��\k}��(S~��_�}�y4e��Ϲ�������qG��@j�͉w-�~��6u��,����g�G]p�����o`H=���m��,P9y��h�Aw�����Q���+��(3��I��c�µ��̹�mX.ر-Y�k��-/K��3�MJT�*��r�>�}���x���øLK��@JTyI]n�[]TS���@�@�Q��a�)��`vo|�>5ǈ�C0:�p�+�wX{���HP9���&����I�~˲l&��,���c��䠀�.t+��Zx�>���q)
j��ǋ����r�N�{1�6
*��OZ��b~44� 2'�}y��N�H��Aη|O��ηO��B���r�ű!��ȰX��4��A ������L��]��<s���ŬH�DW]N��᱿����<4��("d��o��"ޕ0D|�l>�4t��+��ep��������3�RᛘkpI��b�[�a}rn�	ʏ����I'�\]�Dس�t��<�/W'�����k�aV>���\�8��yK�f��0�V���� ��T#����SO3�N8*�d�[7���[�&3�/��QO�����'�e����2����Q�$��@�H��o�Ò=i֢�c8MЇ<�rh�m�ڥ���