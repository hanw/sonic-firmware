��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z��!�4����IE�Dex���!����>��+m���r��yB���sR�~)����MB%x��`-�ȝb"�9Py(>����/{Գ���L�)H�������ŐIыN�����T�7t�Z��cT��0�AY'Cg:Qg�,S�u�s���[OF��1+�}�g�fUea�Ԅ��uPE7a$��n8w�95[̄������iQ�f����7���
�Hr\j���v��~��v��y�A���~|��=/�L1�s�/(pܙ���$�QX^i<�R$@EJ�*�{O�*�C��/�v�z�����5R;��@;L�P��s���wW��=K�¶��s�U��h������#� ���mD �$WD�%�;DB+w�1u���Vޝ܈��e��~� <4���N��I~o.����j�� \����I�6���U�[�����t�+v�g�ɴ����r#$%��@��'XY��\���#S�nכ�[���-�GY[LJF,Fn9�82!��L�r:O#H����V{��Kz��"�@|~�8[��*M�R�b
M�u*�2sA?��~b��ʩo(�EnFS$��N򷒚��W����D���2�:ka6�',d�x��c�MF��\=���q_���etm\:�S�9��K|? ��4Ԇ�όCC��'��C��.��T�l]�īP&K�x"*���sq�%d��47J�k�4�&�Q.{���v
�����������3�:2��Ѣ)r?�z�������G ��z���JgZ�ث)d�@m�����U�tX嘠H)M\�p5�9"E�jK����)7��o�M��+�;�5�i�L���G��)&���_��Z��/�j��WE�N�� �hf=�o^��C�4��eK�ӛQ��0:-���'�@9�K�^B�NX	�	n�uCmY�!�S��vQ�i��/�Z��{���u�Q� �7�1�|��g��U��?Mw�БKC��pL��/������}�C7�����>p��kh�(��K+���#{�s���}	K�e�/p���(3<���𐬜��М�=�ӈ]r��-9NY�����6��'3@��]��������%HJ\����yi��h�Bk&lX|E��xh�}By~�W�ݫ� �� `�KUZ��dS��-,�GGV��m���;���C��im�Z�t4s���YA=h�(��X����U3�]�iE�׶6�7���y�a�3�)���trzX����&Nˮ�����T���}7ʆ��ň%?'�v�	���f�;HaƋ����Z���X���p]��6`r*���K}�6 _����A�$��I���&��) �q�וЋ72�&a\թ~� �T3�#��v
�	��-�ï��]ٖ/O�����skjYl۴����yW;��>�x���+[|Y!]�5��	W@����j�ȋ^���w�LXǄ�X-�Z5�%�-�yv��R�$�����y�d���"|zU'F�ٓ��0G�T�*vn���R43/u��C"3��eWx��;����{�'=���Z��2�Kգ��͝j��N�	��l~"��OCj�A�voP���$�1p�^���T+u�l�#�������t�9J�Ѩ��]�I�T���Us�!�X|���s�ƴ�����
�>ڳ��nX:4�&�-=����B)q�$��%��Y��� ���.�+�?'+949i$O��X�y����տ
^�y�$�섈�m/xV`Qe��@����[Qw`hw����D��9����Rc�6O�e�4��4&�����<�!�4����#B	]�Y/�*?c��N�,�;c-�{Jx���Tӌ�݌1���p�YHo:������oX����4�r��	��vo� �n���?6�1�NR�oe���@��(��.�W��1�q~Ғ���,������ ����$�RO�D�9�og�l8�����mqÔm5b���V�l�x.��`�d/�Dr��q)�����3LJh��q7�>��z�vi>lXt���ՠ#��|R;��dd�U���C�j=U��D�n)�X��F-��L�k�q��蝌N�+d���z�P[�9$W�� 5�ĆSPҚf}o����t�2Nq�U���FC��v����~��c�����cz@�b�9��?���XS�q	 �Ӗ�������)��3��7B�5}r/Q�������H���3���;_p��H-��Q���ڿ���i��5Ud�y�r����� C+o������NR�?d1�i�+!�^�Vv�͔Ͳ��D>�c�H<��3��?���lf��0����tR�z��HD�E7{0�����\]���Ev��:�D?+]�P���dn�����XW�����v	�n�q������<��l������%�Ԅ?��p��fj�W���Сĕl�9���f�'����AX ���ڗ��κ{*�B�࢕B7�t���㻌�¾	)��Vw㰛I��p�.���x�o,��X\�;v�����(ϻ>X��c��,B�k�Zp���T<�.\�-��-ьe�N�RS]{����^�h�����*�?A�dm��\3��HO�LB��]�־�H��).kW�Z?t-G�}v�G�.NV$U ���.v�����������/Te�h�d�O�9��)Ɔ3�t������DhK����Z7�\��ޅ��m��o�k��7���u$�L[��m3�����Pꆠ����b_m����r��/��sm��h����;3�W���m��[G&�lM1��^,��9ɽ^`�h;$��/��c�jg
o��Z_E/�ìp=�0a�<�UE��	�]R(��U}¯������b=7�\-(?��i0�G��`"S���EDGM�٥��)�8�,��(������I���؂��U������G��M�1���2p���,1+����'����RH�ɎB?��?��gg�	�6�w���^�f��n,�ݍ����ɮ�L�j���~�Z���V��G���%י���A_76��5N���2u�cc�AU��`�C�j�U" a�)�
���ζ�2���3��w��� -ף9��ص�h��g󵜒C 쾢�%�0�`@�J{�ݳ`Ei�-�0~��I��mV��u��!,~�R�P�6��-'cY�Ep����|��M�3)� +)~�$\І��#E���sWٖ��s����^-
�nkަ�1�!9���7��$R ¢�����.m%&V��'6�_B��1G:s��뱂nc�dd��y���
�`�R.��P��]�$���D|��=��'\�����Fy&Qs��z�
Pј'
2�Ibw�plѱ ��*}�5Z�e)������8�.�g��+rR�	�$B1M��:Z˹xI�T�/�C}zj�>��5"�o�sJ��C�w����M�m�*|�Ӥ)l�Y��ƒ���%6ֈ
�����n��C"��}-X]��U��ϭw�,;��)ϴ����٘r�Cx�S+V��̕>�+_ ��cg���Q�-�WWF����Q=����fo��:V��RT^|󚩽y`kg݋�ݜ�]S@��3 Jc�q[f!�Y�g�3��#F��X�����Ԫ<���H2�����D��,��&�A���Ӕ�E�A,0����-nR��,Ï�G�bDZD���B*�� �(�ܱ�0�S�pp�98,f���jӤ����^@dNg7�q�3���֬ؓM�v�:�
e��?�
���{m�]�>�W��2yd���*ь�;�c+� �Or�#��5Z�T u��\G�5О&6�qoŘ.R�mt�4���䤡��'R@&w۲���E�ʭ�TUi���Q2&?>��T	��͂Mm�{��eثo2��Cw(���6�ԅ!�m�6�j�lF=F|����/�O�
lD.T.�pi!q��-��y����Fs'�{��~a�p�YrUy���Q����%5�&�6�u��V����uʛ���K��A¶����i�G���9Y�-�,����#xs._��u�D� �G|(�E*�6-�c��#xPp(����6��hБ.��)uQ�����n{:M;6�ե0��mC���K�)�n��-��,A�I)i��Q�L�vVz�L@s�0Y�!��4�7����y��I����K�،��ƛMV�T�w�K�Slɭ뜙�!#k�~�_�%�rŎ+K�lDw�n�$�L�Zg3����q�L�R)񖢕�p:�1�6ra����B�r�Jh�P&D�=5C����4�O���賆��?�Z%k��P�k'*�{5c���K�����~�k�s���s���zr���3�o��F1�%B�F'%jfU����	�&�9�X�� ���3�k��1���pM�+N�}A�f���A2�^w-t{	Zxo�	Z�	�o�U�68nT���^޿2ƿ l{ͥ���\�D@&�"�n���H^��(ᦐ��}M::�t�1�������F\s�]*R��H�Q ��3T�������ե�����ų"�k:���w饚���3�R+�LO�$9�-�>lB�c��a㊌���3�$Ǩ=��#�H�D�����N �]	
�yZ�N�� �FZ�VM�n$�XȐ�Wmi�ᬎ�		N3�AD�Ĕ�4��ʂ+����Q��Rչ
Oǀ��kO���+3���<5Jϼ�	�8��d^�Eה��*��nU�7�'����Oƕ4lb�RU>��7##<)
��[9!c	��b�U�:Txҫ���� Y�v`5�̪�^Btl:;�e�=J�d<��>���K�JN%gi}a	'���+��J���O�g�lC9�d��o��m�����WG[�&���F�	�-�afM��|�M����b��D/�Fg]vX����;XP���o&gK�֩gc�.���	^��Y�Ad���+W�~%��K�;ً�kou�2�j�=r�I�|o�V�F-Hڕ�����1^,XW*3��H)�nY�G��o˶g:�X��D:���Eޏ���yE=���^��UIq����F{�Gm���R[d]K���p������h��V�*KEſ�,��=�^�ƥ{I��Jj�.�[�H��H�Ҩ�;��V|n���&͵`�d��c��>�)2���Q[���^B���Eڄ���P�%R�V�g�����w��!�O���J�_�q__�q������n��o���%�6�F����r�zK����y��;A��k��q����Y��S�w<7F@>q��9,C�6�V微cE(.8T���m�㰪�����Z��@c$����˪Dgn�����ޚ����c{���۳�zV�hv?���`�E�Jٶ]+@��/p������jR��$�0xYί=�����"Ye�ԧ2�K��^n\��gT/"��Iٛf�������a�ӗ������ ^5���CK�gҘ1�ၹ�0.U�����	m3�wU�;��2�.�|�۷=(�)��d�F�l��RN!4gM��Jr��ևKJ�j�����$����}Қ�-�3���!�K�g�Ni�v-gn^D�HR�m��w�)��P�	;F�g�Ld�#q(0��ﶢ2O�>����O�@eiq�n�8�	|�{��E�Rˏ�v���ϦV坰]�U����s�;Wڷ����\��OiPZ�L!���ݸW5�e��um"�!?��t�����n��6�ӿ���zȨ{!L�+������8�$����ȭE���a��R){���m_	�֏�����d��N5W�C5iU���mV�п�cԩ��3�@fn��k#4�G ''V;����	O!	�m�C��[�
��Վ���>o�iѹE�k4r�_�(�LѺt#)ZqW?~����5b��w�Y���z���o4��K�v�_7��DO[%�f9�����b��'૿������p}� 5��뭮&&1�k����k��9��i����T������d�6��fy��p�0ɏ�Dzrzjܓ��Xlu��RJ��}��{r3J�
��<Z~�N��RT�ʯ��8rU�Wa�׆y�AGh=oج�G#x������?�]�O)�"J�uQ�bH�;]_��S��B�	���]��/��=�[sY�����&ߝ�R�{�C��e�L#����uj��S]?#��9Ɂ|�iWZ6;����q��d�ww	 ��W�Kߟ�}�6q�+d@q7� x��9�����~*�uG��Z���Ιh���Ho3AvNn��r��Ot.x�@8Su�>�K��