��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z��K���v���|w���X�SZ2��`���m��o0������Xz�f�Ɗ�P4[i�~|˰k�='1*�K�r�ƅ����o
�r$&���M�/�Z�Lf)��\l���Ο[@v�u`�17�5�T(z�����GI��G�Ճ�JC��}4%b�t����0�ΪM��0Gc4��w��㋫��v?RtU��w�/4�Ҟ��5���wS�bQ�]�;���8�>��]3#�Z����J�����s�\�\~q�0�{�(�/���W~�0f��E��=	
�`䪪���B�m��a�B'���i�S��a��(&�����3>�� 5SB�Bwp�ʖ[��3@S/�Z��t��QoF���b�0i5��� �L�L$���o[��e�1̱5Y�!�D!!�����h+R
@�w����Y`Z֡��I�S�_�S��R��"}z}��D�/D8C�l���M���p(�V���W'�����Ë����A��?�:�u2��s�I��%��-�I}&�1[Sg䊑�:6����rQ.� �b�Y�DH���F_J�`��D�FLJTLaF�����O�0�,ԴDW�z���<YN���EKΔ(�&��D�v�kq>�	��e��֭��8gS�	a�}�障�e����������a+�&�&�: 7ʊ�IA �fU��(Š{����x���b������%�r4v���j(�$�����N�Z{Hm��0s:�^u�ٰcDdDV��u�<�T1X�?e�zp��>�*�ښ6�V2+��&g�־I��@-f7e��=ʯ2s�>r�{ �[�����Si�n³?�U\+�o͂T�W��b�o�6o�O :�=B	V��.n���MLI��bQ�
I=�ܖ0�d�Ky\c.�n%0SOt�&��)����v؋\V^o%� b�7�=�H��m�V��ڄjY�QZ�� z ���Z(�~#)�Q0RY9L�`��ZZ���✴� �S}��7��q�LP����bg��Tw{�a��x���KZ���"�;�2�r���fH �v���"���-���/��Nf$�ޣ���������NsM(���%��)svp�I��<��{��O-j�1K:#�xm�=�J[��Ƕ0���1BJЗ������5ܒ|�u��u��T�%�%U��I$v-ٞS���)����K��j<�We��|��N��O��=�Ah��D�V|���ψ�=�2���JG�;8%"gC��>73/T�nM��0�`�y�̢����ߍK�}sW1!'��l)2�'��� ��n6V�v��/Z>P�L:i����T\: {y�'m�B���f���n嶯!�p<Y��nz-rW����9�nAߦj��dRM왖.	��l)4�Y�+g��m�6����@�9
�j�OO�k�v���K��>Kؘ)ڐK��G7O�_��qX��Rp����W��J�ٓ7���Q�N�Σ��k�w�u�0#���"����?���`�239�����z�`��M�.�D=L`���,&�}x�)T�ԟ��6�w�CI�[��Ѓ���4�$Y�^nkK����جx���Y>���R]�)悄����2�ǊY� ���ח�Lt�j���T���,��Z=_���2�~�V&�5�`����0_���bT���Y�|L�t#0�}�'k�m���͞��f�'��2|el�%�.�G�d�]m���Kr�Uޘ1�R��c���jf���������0�1��v�-��
l�r�2�$dh�I��ig��.o%j�q4���Aq�2��g�Hw�]`�}N���Oa��ݎ�CV�����Q� ��]�X������ʲFD�(]�W&�,�<�Ws�g��ۂ���i�FA$4�l����_�|o��`�ף����������{I�Z~��sO��m^����<�׫���W/�c�;Kz�h��f���y�j�&j��[ȑ�u���Ҳ��Xe�]h;����AgA�z�Zx�e�@\4;)�!��D��=X �֨j��X0�;�'b�/�p[�V49�c����Piny~K�ꏖ�ꏀF^^~_h6�#��p!��T�=�%'�i�ī��vr	��i�Κ�4 8BÀ_�r��ٳA��뷃Nqb���9�i� y�����?�����R��yJ
I�L�O��T�>J�zr@->/�����űg�rNG9�$D���d�>T<K{\��7���q��ʃZ=���ֆ�'��-����9���Ł���B�2����ȯ)6�k��`��o�A*�Y�Iڨ�<D���x{7=q?T­�,B�} f�9>m(�0�?��Ȭ�|H��SBy���h����('��xd;Z09r�}�O>*�	��R�]0P7�A�S0�@�|}T�`w*K�P��ȧ`7�bv�3i�{�#y
(�q}0�G�����&ӝ�k�?h�,�����B%�N��SX��{��]4�z����w�Yu�|ҋ\���\K��Aɦu�zƔY��(�A�@l" ��^¨j@'x����g��֔F�#���~q�\-��\��6������zB�$"ba�e�-`��*rT���7ڍ�T�x�KOs���G2�~hc��7�w��Rԟ����iw!i+��Dz�o夤������ڄ-R�	����#�b�eߑR���c��8��Z��W`�\l�hl�Ƥ�B7Q6�/!�:+<�=o���|���8:ꡑ�IRwT��'�M2K2�:��.�k�@�'������mR��C��è�C��#�����~u%��_	�H`����ڔ�J+Q�W��c�v��6C״wW�B�Kpm���4}Ry)�1-V���r�bfǤ�y�7X/�A�˲� �Z�6;���'��5.� ��}!��vo����|��g����l{��N�i/�w�6���*�GM6�<��k��I�;�����&?��FyCF 3���o�l��l�D��N��i��v��Ð�6?a(����HL\�K�_(�63�-���0� ��t��$}ݖ)I����9���j���V�.:A^j��jfi[��E���#�l��}EW�@��}���"�#�1��F��"���j.I�r����N���ߞ�=���觲7)�=?�"*/��B.�� ���&��sR�oEQX�*�SRSC2�%�lh�����5u�8���~&^�a�s|��)��Go��8�e趤��D�k�	������o��i�|�m��«��i�Y����}7 \�����F�|~DX�O�-X��'4��D�7�/��c�j���݊���D�y��]�0AU�DCG�)D>o9wLl`~<!�z� H�O�����&@�;Gjz7az'$��
�(ϒ���Ӏ�B��ϝƊ�K��ɟT���������,C�QK� 2��mq�u�z�F�����@�u5S��j&�ڻ���K[b�'�*�d����~W5{���@P��V��7�/�\ݤ��}�%N�C�M�� �\�?.9�L�9@�Xh)�����ϛ�1i�޶ى���)������"  p�	ZCk��Q�����Asۉ��Ł�u��%����Ȓ:���U߭��ǅTH�ʹy�y��\�EUUa�ss�{}��Ym�6	�e�<�DZ %Q��¡�0�ъ�X9��Yð�qE��!��ɶ��MP��k�k2�=�6��L�g�� !�q��#�2���us`z����������̧�sʽ .�:i�r>k2hJa�3�^��~������ۦ�D���K��>g^־!!)�`[�t'-���8�(���<e�G^�	9I��̚q���;�Eq�R�y�;s��9M���&�`^kZ�
w�	�<��XT��SF��E�����q�7�l���Gw��0��)��ac�3y�?�/�X�A�c;�Դ|I�J��\�M��W����/G�Z��z���?�T�d��!�\LZ����gׂ\�he�)P�o���v5Nǋj���;W��.7��Jc��쯦5�';\�d_4{J�z���U�7VI}g5Q�!H��H����.dB�w��U�^b�4�Ba�]]��4lG��ݿ�!ß�ټX�~�K���6\��W�n��S�&1�P�/Y�-v��M�s��L�c��+!O�r%��=f�w\���k�<��RKݤ��Z'>Tۈ:w�{�R^�Uc�h���K�ss�Aw˩R�@i���>&k^g^��9 ˳O�������zG����Y�,��J��̨iRa��^���&ןr�ᅫ��<$��(}(�tZ}����b_����ڦ�HC[�A��`1;`<�0��>yj�����
G�y��HjC� �?��mM$��F��eڨF�Y���$���U�4��u�F��wEG	I-�ga-��A����/�g� �u4m��W�A�H	�^;l^�q
�7�VR�=� ��}G�U�)���(\XpNn���,��硨9�\W�?T�Qq�-�@�Ğ��6�����M��f�>(RD|Z��5�)���«o�J<�f�-��Jf�R�e+=��6s��^��tz��'[)�8=��k��n�F�$5��T�جzyY4[h��-u�E8"�gk��G�<��wj���q7���F阇��k|1,
/�e�D5���O�cI?C����7E&9�֝_�(ZɄ)t�8��Zl�"��>n�� fܫ8�Ɛ�k�ɐ��tڨU� �&NZ�%J,HvQ��E���̓��N����<֥���]�o�+�����4��w�3���8���	���+-R"��g·��9�xJ��񆮉/	��H	AR d��`8��vjxU�)��:��n�̮|�(=�5dax�f���b�i#���^� � ��Z]�5RW&�忛�+�K��=�~E��I�}l��B��WꋉXʗ���t�� �����Qy)�H����v��E�f�L����V�^�H_Qj��;J#��28�P�p�Ì�k?m�܀���F�@*����AvԏY»�������5���e���P �*�TQE��9a݃]�7.^Dr�y{Or�a=ņt��y�Z3�Z��xg��M�Z�>�#vF����x�a��_~�\�LKM��nF�פ���34ʲ�岾���}ci���0k�6���"�%��i�����>�?}u�A�oZů1�nflQ5�ԀXI+���#0�4v��#}�FW^T�nl�$�*O�s �f)7�WT%��Y�<�C  ?외�|ej��A������y���e�i�@eQS@�$� [[͒;�D%=BW��c�CW�r�����5Ef���ֵ����j�@��
��F��RT��7c/��q (C�Vp �H�/��2�TC���`̗�P�A��q*�R�8ѷH+�Zln�_I�@��F�
Z$Z�y�㴛���k��lU�k��4#ֶ���J�k�$=u��.��L�1lQT�Zw�c�U��Z(���f�mr��x��O��`.4�f{��a���P��@�*�:���J�z�~?M�H��x`��iO�~�F�=��Z�ޮ2�G���H���>�R$��<o��I����׈ô&��;Ņ���ߌ|Uk���7���*�X1
��
0\��Y
x}$���wٳA����o���v���$� g�,}L��˓���Q����eiT�]X��5�S����L�!Mê�x]�`��E��M!H&�|�6���8��K� ��� V�5"~c���AO	�65���]ow��:y�6�}���?ꜿ����]b�A���Əu��{�u�I�<�<D�8��{#�rD%?��<z1�S +�$y��>����*�ut}�����\��Y�o��T���ξ9����!�c���Ӻ�>U���+qĹ#l�o�W�7����A�*}�`�L�* {z�����7���k�G�,U���J sM>99��3����[��`�l��Ù���_1\5t��C'Lt!^�6N P�*�Y,�S�C6-���c���V�b@/,�����n��*���_�9�u��2�s��ٗ��"|�>�C�Q��a�L��>�2ݜ���E�$sZ +�)\3v�.+�����?ξ�����y���(�y@����z�[���.���?3�?����p�ߏ�"꙱�va�L1�]�Vr�B���`mC��������.U=")����A<��@T��I��ij������z�k�{ʄ�A�p8���o�f�T�&�T�ё�vI��n�y.��%cs�+J� B@���'�uKy�R$�
4���zɥ�t�����>�Zѫ�Y��yN{� QAN	C>҃�}Z���9�L�dm��/b�`���gmUC�hiTp�����>�������6Ȉ!�Y����!�H�y�i�(��\�]�����.�n��SCE�9�&ֿ��"��(�J�|�'��܀6�A܊��ƣ�Y�b���ω��	����b��H2�� v?�?�s��5�/%I�DMqG�
�]G�J���5�բ!@Vjkni��J�9�K��4Mp�ƙhf��O]Di>� j�|�����*�rt��T�N�ϒ3�.`�G4��bT�����F:�E(�;�"�9f�s��$����hy�H���5�.&�fd~D+�W}W0t���{N�O����Z�VE�1�7F+k�iv�$V��ww �y�D��{��"��7]��i%4���6�w�]�А���%w�c�P�-8��b��h��*��}
.��Ͳ�1	�D����b�O�@�w�1��P1h�Zo��;�y1MtS��Q�����Ic3�*h�:�(��� �������R��\b��96>��R� KR�z�lI���n�uo�ZK�Ar.�
9?�̋����;O��^�LzXJ��ժ���ൊYD�:g!po�ƽ�M����<��Ƞ�l��/4	�!{ࢻFG�O�������B��/0��Աq�0&q`�f��~h�ٿ&��Ht� o,A.�i���O��aB;2		\^����Q��~�����}�j��^�0ɖ�n*Y���T��q\H����dk��-^��ap"�������w��-.	��wKI��e7�����U_�M4q�KS&s�H��W��7�����nw��K9�_5�7m3��6|&�S�����YS��	�,�g�a/@�����W��"wR����~y��C^���W_<��F�4^*6��+��'�J;�B����G(�W��iXgb5]j&���t��-&��p��S���+���Z�|�@-m�W�.�(>Cґ� CϦO9��lacfH=�ʞc�3� %��Æ��U.Ϣ\�}�$��͹_��*�g�Ӓ��T:)W�Ҡ��:j�ϟ���e��Y<S��.��@���=h[[`�
#U���:8���i�~W4�_V-���5��
�>J���+=�O����?���I�Z���>��8�� �c�B�h���VG�Z���y���!�&`Xƣ�t@3u�F�o�@/�٩΄������Y����g�*�в�\@�F[)儢j�=CMܪ$�\���D1v �FpfP�_>
�v�WF��"�ί2��u��;��A��+�3�.�E�F�s�����g�V�z�h�����	5w��W[�����e?[~�tgM*q�{/e�o�'ϛM�PN���P� e�k2�1*��y:S�� �A�^��	̚.��,����7�P�}6+?;_�3��{*�9��Ռ�c
���;�Z�q�7��+*�Vt������KN | ��q������m/�ЄG]8�#EZ"����"��:Uq�82[&F���DiY�on�9��:�J��0��A���I
S�|Y#E��+H���i�E	w ���$���ְ߾K2�
�������h}EP���x#+%��kX�X�Fu���H)pe�IGii�E�pj��&��J�Ģ�P�Uh(^e���|x��@4� ���' #�>�l];�g��ש!"�Z���z��f�Ø��UP�R�=�����6d��J��@ |�R��O��� ^B�V�E.������̱�RES2ԙ�=�K��~ϳ2c�����qeD	á�~t��0��Z�L�
��[		�E}U+zͫ�,ك̵���'d՜U�8ج�Ǡ��7�,K�!'A�������+�3�ȿ���K'V��b`rIZ�v�܏����t��coC����P��qf�=�_�&�����~b5EqS��(�p��!�G\�����XS]?�!X������{Y���c���׾+�&�aÚ�7�	=*u&X�{.�����L�w����Z3Ԕ	��*DE�^�۹��|�"9��}u��2K�5�E[J1��z�Zު3P1�� 	>2��9����sJ���K�BQ����EʄT�2�QB8�,�����۷�:��w��k�viSg���x�M���$J�$zaT��Vf��|lMj�=�R[��w� �A�c�gY��A)��'9ޘz�-�N�K��зC6ߒ���ǁ���C�lB�"*��ciޢ��� 쌳�4sү���(FC>"�2�6�m��<=�Mp�O�)���a~��
Z��l�m�h��9t��.�N5�jf����39����֖�lm���w	4�!'�����!~��(���}�+�D�� �p������1W�+�^�(�N}���`��̹��hVDjU�}0����Hn�H���Cdd9naް��6q��$�lF�Ά�������Ц��$Z������se5�X����B���,���83^^	RRH���_��>C�����sOW� Fǿ���P��5��^Q��QX������r��7�v��	�M�r57�7/����2ш׼^��d�P��R�gOK�kҕ��(k�Շ4|�6��Ts�!U-�����<�hq��0ٸq������QGHg��Z��~��Ș�:��-�B����D[�N��@;0I�X�	��E�_�u���l;��K>šm_�X���#:�# }�;�lWH�����*M���`v���-4��wN�R�Kf|n]5�����_�$3(<��ϟu�V?j�� #.$ng5��y �6aP��_̈n=^ʐ�vʻ�F�[&n��v���9�؈�q͝��$���<��4��Ivv꼼j�b�&�b@?'����<�jQ�ZhpMH8eɤ��$�Q#Pϴ�����|�� ����gy�E���Z�����e�(�fA�ߩ�k2^[&$������W��/�2@�{)�� ��RfjZrn��c'�u[�3�{}Fsm��	�y�������]$!�.�@-/��p��x��e�ռD?�ؠo.�Y�M!{H/��`���ό<�^�g�fn}?HV|*�23.iƵ��o<�T���}/�ڍJ�͎�^����1E��N�llyc��Llۋn�x��Y����R��s�B����L���3�Xo�0`}�J�O��3��]��9���U8H�^�����8�%
CY��:���:��{���m���~�8����\Ԯ\k1����l������xfT�#r5,�y�-����lc^�&#���&�;�ș�X���wTp�݌[OQ��^OoX�e��/��l�Fw\����J�f����.�)B�.�Ř���p�����V��{ �Ƚ�q���u�&�Oji�%\��[��`Ng��}�\��y�ϒ6���#�fv'IFdGE��}���ݽB���z���m]��+?�q�&�I�!SP4��Y�X��CR?�F�na�庉�c�Ȭ�C/��؀lҺ�ʻ�,�x[9��E@$�&h�������J�<�$�~��(p��*dIw�0)"�I��Y d_�&u�
Ƃk����.�s,bL�8�k㷶֛���b�+7g	9�\��:8d;���N�!���!�M���+H�����Y���|zhjY��#Sd�'��)���߹[��,���s�a��×����y��ի�����3��Q��*�ߛ#L����w�U�oŷG���/�n-d�w� I ��**�2d��4~C�
Z��I���ȷ�,�1���䫅�`aB�Q����C�/���Ab����SU&ڷ���ST�ZӺ���%$�f��h��-GN��(����(E��8H�ԝ�$Z2_Y�����F���i��~�qފ�^q|��~m�Pq�~�]��؝.��*C�O
�	�}	l�*�Ds����R�Od5ƂrT� ���(�#��iIpV4l�8E&��& �����/	�N�B!Z'2��"�c8��Jjs��w�/i�	`w���<�Rah�.�S[8��Q�8*���lK�����+�[B3��Ok:���ֱs�=�o���x\�T�焮^@��!�-�$�E���:+�����a�|���*�(�&��!8E�(�Ԉ�a���C�iUu@Y��5o��e=�q�c���K:H���\ןr�S�B�n8�~qui�Z�Ak���bl5g��zH�y�r2UR�1�Mll��w��'8�!�ɅO�S�UD�uc��(��b�[q���罸h�U��'�1�{X�j�p�.�Gqk�~��F5VFes��n��7þ�:�hjg�Lfڽ�z7�
�U�S$
]c/�T�l�7��H�bT�yc��Ae��1QE�����0������n0����yjv>�m6�$�?��N��[(�&�Y�x�TV���&ti-����\������	�Ѡ �{ژ�~IcvO��;��B⫇��8ֻ�F����&H�X�I��������Jy)³��J�iQ9u��qz�m���������L��K�܀�$D��A&>m�c��U�(���E�]�.Q8Om�"|}�;{ht�`�QJ2���e� ���W�.h�_��9d����x�~Fge� >�G+i#���q�s�q���#���he�O`VbJ�Nm�;B��'!���K�ߒ��H֝D��'����s�]��rT�$�u���c����e�8��ժFs}n��_&��C�*�d���Q��j81��m-���x�`X��Io�;�f���c_���!ԏ�mDV�u݃�?�(�n�����Ț%�%��G��%+̐E矉�s�g@�!�HD�����C��f�t�õg��\���u��@� �/�YB�e�S��'�F�)�9ֹyD?+���-���B����f�뱌M�U����'��)�c�͋0۬R;�:��҇b��{��XJs3O�$�3����c�!�Ͳ>���-����/6D$͆
�����K/[m�5`,ʪF7%#��ƈu�lGi`Mb��8c��6$s Zw��y���pm�NY;�f�h]����a}O���Ҕ������E=!냪�6\�^'�|�{��S����?fGw�4��s��U���וp�����-⦥z�`nNr.R}<5K�����������7��z�����]u�sӴ��d�$�o�)�;�d��_�NPxɠ�Rl;�i�Vճ�� ��s��/��dz�fO���%.RQ�.u�ޜy���O�j~}�11�	�\���b�����/�/Z̨NE��cz�-s=����O�W��?B ��JW6ĔE��ؔ�����{�zp���Чb��d[f�e���#�U�[�"�N��5{lϜI݇���.z�R�B{�6r0��N�6A
���N�\&����*	����\N��:(�?% ���-��R�c��ɓM���m��0��`�(>#�3�"	�x	y���2-�d/a"����,ZDe���+]3���K�
���.�Ye�M�ο/FӞd/��
���q&��V*8ޒ*U҄��Ѡۧ�w��v�&�54����tr�#;J[��v��tr�bb�i�m��rѩ�6�S�M}�5ٿ��<��lH�=���T�7�?����<#A�
�;?��ٖ0+�o��&�KP,�ba6�Am���T����޳�Á�C��Cb�(	�ɨ)���X~���R�5��XW1�P?8��Esi��0}_WP���m������-�Z���_��w� ;��/����Q6��ܗ������[�G��[�0ND|�ˉ�/���1��ʉ�*p~n:����skEB��&Q��B$#�6D�<4[���Z�3Xe���22�~"��:����S�tp�5��|�\Y
���w�ܮ'>1�r�x=V��m�'p���P߄�Y���0ґs��ǧ�W���@��_V6څ�jPݞ�;�X��Y��m��xq#պ��q�[��T��RF�2D�2��U�l�%�Y��o�_ZGM��uU3�E@sCA��{G>+���%�
��	����٬DP�R*u��=X�+<R2�%�\�t�Llq�=z0-�A�����L����b������F����b�%��#�'�],
�QH0��Am>.�у(���t�%�
GW�d����AA����O�,�/����'�`�1���Yj�����G��O"�7��0FG�q��!��mOiT���u�%}q~DP����8�%�J�~9#��L0��$���Ox����bH1�Z�C��^�h�����h�qT��I���e�٨b�E\&�b9e9Ӌ�D+�B�Z���9�/{�b@�����\W�D9X�z7�ʿ"1�ss�XM�g����T5�#��|M^�fh��UE3�2��� ����N�3Hr������D<�ҝ����:I�@��ȪhHS�ґVs��Q��YȤc���X���T[�d7P��z��#"%�Pf+ZDQ�\������O5����i�O��l%&h�I���y��(�X�� ��N)��%���Ԣ�9�0$�Q�/�C�P�����w��9<���A��,ѫ>�E7��s||�@���csɩDz���V��S��ђ*��W��rMh� E+�7{�Կ����.N8�J�[�n��g���4����1����3�:��Fʐj*a�_yu�	���J�n�,N���<���*���J:;.�	����P-��|�FI��3����w�!��D�W�]��􆪳3�ZX��/����(�E/n=3Zr�ĕ;>�g�⦫�s�	�����3Ѻ9A������8���")wr֮/}ma8g�����ŏ�=񫉳�s���Y��@�Lr-��mz��Ր~M �e .�W�~_����>^��E�VZ�1���|uj|K@Imtb�Z�>����1�y�г��F!����!�e�W�K!"`�_:�v�`�������ފ�7��p7��K���I��N��?��v�G�Nۯ�����/�`5]ϧ��K��lΌ�r�k��BR1��J�0l}vME�yP/z��[��
+���Q@&0'�f��:�=��Z	�8��W\��*,'�%l%Ǯ�<ɗRI�=��O>W7Ys<eP�D��w��f~H �!h�˜m��Q� �}p�ZݓyO?ǃ�� `�U	ھ�]���4�V�(F(���܄*� �_]��p�0��Mn�C�ٲ[ӕ��g�K+�P;(�:S�
M]�xF�%�W�ߎgBB�QP��(7�%2n�ߞ��iaU�Zb؈��/�D�b�����6#����RyKF��^"��G��B;��h���n�v����2�:iA�����^� Z
��47�V7����l-�d}���pA8�i��$��C�ȕɅ�xV�T�'LTd��X�T!'Yu�/��}�5���ì�Fb�+�P�����*sy���٠��H|4t����ĥ!|�(ݣ�h�,���ͲJ�~���:~Z�dN���:�(ם���(T�A������q���3���{���\!���Q��K{J��)®؜Z?�ď&�
`�bg�^�LUM��w�J��dՉ�H�Ԫ�>�v ᘸ\�.'��m�_v<���b�
��~�F�A���ʙ������%D��7}�I����&a-����6`�*�*b�\�^����\����xy�DN=1�E�oo$����7F�ґAw��/nEQrH�݁
u�-�W����Zv �
+��ǈ�3�������g��hGR��b7�f�Dz�iȡ7\2�x�Zځ:����n�E\��c��L�y��r��u���2(�����{_rq�����8{�S��Y�ųI�8��3]q�R^&_V�^|M�e���/�[=BLW�a$�G�D����l/�y-C
��g�s�~�0�w$��a�гݎM�V���
�@w�y\���vtE�I��.����!���s�*���$��MY���F��w��p~�b�|I�n̔奲�ӯ@߬!=ht�!����S%��6
��f<?�,��6���0�660������)+l�ؑ���f�����x�!ߠb~r���U�Ƽb�UN�"	�B̺2� <9�5Ғ��if7�ev#
E�Zx�����z��Q̟垳���PZ��4"h���j�[Y���Ƶ	�#inI����E=9���̩�[
*�H?�/$�[�oŵR�_Tm��%>=� �"�o�Ky��P��N���x�;RW6������	!�����!D:.� ����\���͞�J���+a��e/|���A��i���g"�������1UAp�s@ރ+^�B�����P�G}^>ƊeP��
KP*����-���C������Z�Ŧ] ��������[0ꎅ}f_R��ɧ���Iܘ����/u���k�'@��&�'fJ�[*�ê�v�;����1�i"�`@Nc��E�������sw�X^L��"��\�j���j�FLZ��աN���-��3`E�����)#�h����!�('��V��C�؃�v�nz+2���y�Jn����-@/@�&���2�2��:�{�:������q��Q�\!<h�v��\?���f��4k���fp$�Y�Z'��yo��}�MJK����B���N�o��U���$I�������BB1
�.Y���j.�{b9��m�Y>m����n��o6�G�]�߱�A��u��X"�;��������������D��ΐ#1���}<���O���@{~��|�h�:SI��x����ň����ˌK&�b}3��%���t9�m�>l��n��UkC��:�	]��4%KC,�N��+/-O�zIG�#���I�.��oR[�L���`����� �'�v����/���F`Pz�r�+h��Z�Z�b��>��0Z���]�?�+��s(���톾�PQ�Ժ-r���,q��S6���T�����:���N�/���5uI���ĸ^�b�gEui)��KDs�cDȺ�_=<J����ì�}�]�"2�3���1.U�ߧ��7�=��T�t��L*'������m ���~Xs������\wt���gQ��`���<Q�BU��OgL���'��Wg6�=�� 	����CgU�ɒ�[{Ț=Ւ:�ze�ua��S�.O��>6{"OpcGy)�ĥ�y�@N=�� �����%�?���B�k����������Ү��ZE�4�^H��=��5E�ӁkJ�4�?�?D�4�����z�?���ܮ�&�-��h�\ ��*c(������X�1��?���GMAo�h��3<�������Vؤ_�#b�$�t�"7��y�	j�7dz�_�.	��p�۶Bf(f��A�O�,�ew���
�u�>:��'Ԡ��2ҹ�n�yHL�wQ�B�F%�e}/-'X��hz��Å��`cp��	���7}K�*���E���Մ�[����DS��|�oq��͛�mP��o��B�C�ӕz���F���㟸���c?.:mnj.�Ɂ�;�2 �?��(����%w���g䭂:Q�Ϫn�Wi?Մ
��@ōp]J1,���a��$�4[����U������1<H|&�L����O���';͊PY�o�e�)<�e�JM�Fh����V�:�~���<+��d�o��G�R)82�rN��p(f �T�:��`+8G�p7���u!�ܶ��ND�n@�c�Wf��LMƎv��Sg����`��&�"�{�1�·¹k��N��A|Db~/Oo(��ͽ�E]���	)�2�u��;�� �_�(�S/E�.J����	�W~�i!���#��u����g�D�zN�Y?N�@���0� 0q'@c��8A[p[Gy��!3~P�=	�Ƌbκs�)6����A��m��*�-̻����4��O��ϖ>*j�Q����7{�l�-��FTTJUdSI{7�}��l�0�#yY����PN���"ј`Z_�K����J�N�{�{���o��(RGV�"%�ߚ}~z�i�V�&�p8�Rn�8�m-M����WQA��C��ן��{��I�/����>�=�w$�d�/!�ی&KDBn��V��FǤ��{�U̫q���ntu{HU�r��N!�i�_v;���s��9U��r4܄��[A�mWL]L?�ۅ������:i�L��A�v(t��ʰ�kgL�� Ɛi�F㔎"7.�f!�@^ eQ���x�[��x���!�q��v�T�#윔@2п.�ˢ�:&� =B��RBLtk�)��SƗ�G5�v��7�d.�U`����8L��t��ݦ���O��I	�dbP�+��3U�Ns�Uq:n�q�C��%��R�\���W���~��P����&���*�a��������Ip7Jm���n8��a�Pz�*n],!$��BՙM�2���Jb@��j(�#E��g��s�G3X��P���DWiD��l�A��H�ݠ��WF��Hݺ'1��ؗ�-�q��p�՚5�����N�s�����lGc���}v*�TGh!_����x����of�
�`C��_C������3#�S�[[�Lü�n�v_�,���K�6$�TBB��`��@�@�(�J�,Գ���'���1G�_�����v����9q/��s�A�@Q5bN���n�
-�ML)~��@��R&����)�	b����9�B4��uff��� c����slwqF�Ik ��P0�k;غ���)>�֔���b��^��)�u� !��4E� 꽚�"+(R����ʨ�)�Q��e�P;���G��F.y���	}�"k�#��e�D��q�?��o̳`�X��j$ŒR `�����}|+K����+���@e�����@E+@p��Idz2����Z�bM�`�Z�	W�U
�S	�����k��Oא��T<"J�-���v0�XT�\��mp=n�$oAvC�V����X��~GRp�* �z�ę��m`빇`�����x]��y����k5�>Ǖ����4Z��Y�+1���K�K�V��(�QȢw�����zww��'-W^�CC�F�������M�8�5PQ���>�̝���{���2�`S5C�����`�����>��v9���G�U��#��v�N|�$q0�x	�m)�MG�� r*�6��ԊD�D�G�ֻd5O���*ũ�U�,	6�yGCU �p��W����(j{�l������v}�
����4No�grU"��^րc@�g>�h��K̽*���Xl����L����E�R��3�ڦS���z���=�,H����=(w�\Q9��T���F��l�s_��'�93_6�(�*�(8fϐ3Z�}"J�_����A0���eM5	u��~����ƞ�=M����:�����!�M�E)��"�g⎜��ID8��4��Ghk8����1��G"ע���3ַ�zվo��-�h����{Ԩ_~?��s���i�C!BZL�\yl/Oh�On�1R��r���r0�zs�9����h�N@��2`��驵1q\G�_�D����8
��(D�aOE*#T�8[]�<�}ݗ���.W\�+nsO���E��_奔����(���d�Y���r�0>��:l�u���T,�2���Ɏ��{N���ܜ��Xu����$����#��d��l�&�*�"e�ʮ������I�m�J��{�2�j&U�P�A�x���V0o0Vg�ה>��ٺ:���]�<� h5���,�d�"���)q>H��O⬋����4ɔ��u���Z4߻nsU��ǛE	��7Oȣ&�kW$rJ�rw�x����m��ۨ𙑽K h�-�KW��aG�{���1H9���?jT� �˔�h�7�r�~�EyQ�;t�C��)!��va�<��?i;ʣ�k�?)r�0�L�%,vJ�(r�kO۠q����EQiZ�
�'�va�G���_'#?eK�}F�W�b.�os�m�Ƙ٩�9}V����aju�	$K~�ɖ��bG֌�5��T�3rPmK��S��]��Zޝ̪��:ܨ���S�<Զm����+��=�9��?�"ST�����S�զd�_����}�7�ăm,���'�������?K�?_q	��֠�p���<�ٱy�u�Z(_��L;���eWU���3��W1�n��W"w�}��K[x\z�^�dՅ��"���J�@��q
H�S��j*~�����'Ԉ+V{]ӟ����!��8.�������!$j,`oz��o�r-�\ .H��˙�be��~%6�e�N(�`v�}4��qt�F'AY�}��V-&���z���m�$�>��}?3��c+�a��V���?HF�&��+�<��>�b�O�F[+E���BY
�(����qh(L#R]���q��^<�rQ��0fă\SC���u���.��SS�se-�){�F�E!Qk��G���O��L$�b��65O�#�����+0CL��dG�^��v	!���=D4����2�ң6�0 ��ZN���{���b�7���
�/k��������N� Ä�F��b�\|�@zK]�8�%ewf%CP����f�xb+TL���,�Htb������L�}09�Џ�BHpJ\'y�F/��͒�ثۮe�����{RC}��K:|J�>�Qa�9�{ng�r|����խ���#/��4�E8g�<B���A���o��H�H=�2:��D�ϰ��(��:��z�`�(��'C%��5�=�U]���w�E��������8.�Ety�Z�Q�b����X�r;����ݒt�����$�&�N�0�]��@����r'�#'��{����A~�9��=� �'��
�n��0��܆E^[�}tgwE�ރ�UW�>&�N~4�am�u�b�EI�˘��;��A��V��=�0�0�8�{�Y��� |f���A^	=`���΃6 ;�� ���;*	�Wz�2��s��|��"��U2a��2��:pc��'��6d���ETUJ�ka�Vd�_��j?
�XK��rC_G��m6�� �1��ڦ�u�:�Ϊ�踤I�'��- g��T��z`d9�� f�}�U�8�7Ȑ������DR����K�
��d9��!(i������9sD���TT=���	9h�H�/ͮ.W�B��D����8ϔ���G|�q��&�G���*Ǒo?'�p�S�7 �/%������@ ,^T��v*i���iAY�]^>��0$�Yp�W����;�ť���8%���Ġ�*V"G^�`�צy#��u��)EU-�0��D#��ό�$�J���;�kĘ{vS��6qm����]�; �Y�i]�Z�`�k��ʢ�L[L�q!�>Hm%{u4o�&��9�?-�4�p���b1M;�����
�����E��<_����\�Qʴs�]R;���tp�����	�L]������b./��k	�9W	@S�r:����Ձ��t���U���e{
�5D��qQ����X/G� ʫ<*�!%�N�Fm-�����ݤ>klጀPͱ�r3��;�f��Sa���3�z�T�HK���7��1����,�]���Ԫ��[oZ�HO���I~"��]c�͛f����o�~��v�[��]���X���=2B����=,~�E~K�Æ��Z2�6����B�BB��(R�dq7��nOڀ˂עn���S_jf�g|��ˣ+��w�޶��/���nmz0v]��5j��Df
4�̓uUV*QO�q��Y7�o���L6�\y�1�Q� �S�����7��,���.iZ�<8�l74u�}<�?���D�F�%X�+�J{�K�7Dk��E�C7K���F�,�E��p" m���a��aG��P���\㸨3PQ��Ϧh�wN'k*P����i�KL��AF�B5�W���ل�Q��B;l���!��d]���>ȂY����9m&��	��X�KA7�M��]��&��=I���zj�c�����C��V�
�c�޼P_r�%-�0/��/C�"�Ƀ#�]��'��mL�J�!��b�LG���
�������ߩ�"ɰ�=|�(����9K2��ղ^�@G4=DVBZz.3���c��j,��Ь�?�\eč��_2�"��fLMׄ�9�`.�� G�L?�d��'�U�$��]1��_���
.-�v@�R��%mi~5;�ː�T/���wQm#-����6���ml'ƹ�IA����-P	�P��M�O�OӘO��j��l���B�L��u���;eN�����,�`��=��1�)6e�MI��ȭ%;<B����Ý3����*Se�{
;��$P�7����$�=��(O@K��)�y�V�I��?cN�%�O���^�(�솽�p �x��R�J_� �k �Q��M=��S��x�Y�N+}8]���n���z�����~ϧ�a�EG��{���=کr�)^���`%3W4�޼hSd�좠7�,MC��� xa�.�H���@�H\kXb��(	��&���#;��J���g}�m���*\�W�[�#��WI�K8�4Gi	�ye���_�C�c�y�.A0~����J�T`|�&�J���K#�>���6;f���Z�	˨b4GG3�����INH���IGY��>��PT�J�`+l�х�_8�Ƽ��zh���9�
x�au�F�f��q��C*̵���9��>z�5���~7������gU�y�?[�����,�{���՛hܕ���F�}�Q��eD|��У�п�,cC��\&�{��T�J@�0�	���e�w��cD�r��4I�7�+�ٌ5�	�5%�����(��B�^��0ͩ��I1��@�L��qz����=Ey?;��e��?хbU۸��\B.o٩��h^#_�L��ږ�/�UR8?�d=�uW;幠�$��b�,��H���E�|~?J��X���
�z<�'����fU�
'C�ٚ:R،.K	v�m���{�&�|¡3[N���B�\g�Ե���0�r���"��0dVI����$'1d0��Ӏ�p���G����9����W ����FOI��X
ܖ�o�INふ;6u8J�E3#o��/��-��ݵo{fL 1U�qd�n�� N2f8�H\�,�C�������,9R�3z#�M����t��d��ɱ ��~�Ϧy&f�3m��4x�iRJ����w�b�YGSr=��d��,J��-�uDŴ;F
���Ú(���\k��`*�����apguǿK�԰��%x���H�4?A�4��H�mkR	�7��s4mf�� �>f����5gwG�P��[O:>s���<'~����5h`l��Zc�uF$����$%�Z�F�;��=��6aD<yi([���>��\���_?()��:���\�}k
Z�y=�=t�����<:�ZA�T�<MaJ`�����k���
����T;
6��M���D��V�KY��h�����D?�����(�����N���f���q�M�"�=H0X� D���\W'j��"č׀���������%�Zw�g�|h�B���j$�N�Q��I|C�{ *F7��xj�g�!LQ���!ev/ɲR�R��-�VcE;gl%�H>�5r�����ˑ+~��Z� _��w��,#�	f�$���.�9k��%����蘆��<`�sS�G6"U`��Fh��cYc���-r���f&��1�ё���f�1��P^��_��W�r���PVp̳�_�Yx]�78h�L�3�O�3[�3" 0-$�8_���yk5eO^Ay� �HU��ρ��~nQ��B��E+x��o������$w��wDXxZ���P�XJs�	X!������_��D8����(�1��sk����ў��r��|�����cL�$�B�f����?4�ǭ	��