// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sfD7HCheoadMccpTZvpuKALDzjNCF0Fu0V2yOf5MqH5BvEEnJv8utHk2P0rnURyB
NA/URGvXyHmpv6tfIGXfCrIbFAMTKJDND+aBO22V1jOsTp3WhRHReqzTCknFmIIm
GTCFu01RG+mE25cpTWk0ZO8JqNJkjItfr/7+rC759fo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4544)
ICY7GeodGweldDM8GQzQMAd0yOVEWiXiXgZeASvGocVDTI5RilrGESAmCV4OiDtA
MnJfu1sqSMGX5iC5XHE/2TvQjC3xfz5nuMUa/BPEPzaZyePeEdvjE60eW1I+8u82
rE2zd4YA56pd3357rfkluEhBy37XSdtpWDXMMg8tFyDE+G1X4We43sd6C13BdtUI
pZRvJBBrRinaVGLO+QTgoWj2zFSxfH1cqE41KPdaGE80vNqsglmov5YLLDGaP9/K
5ocLNJ1sRtM8wMZXsUG7BqT/I9f5BHTXsU/AWl2pOVcoNXEwfY3IODOzv+8tVJ82
Yvj6HC1tm8y6p9yfw3pNnI9XfUux4XlU/XwfWkStfxr0pOFRev7fAjmhTPBpqCVa
JnHuOFcNJe1XAehvfL78OOpH4ZpHk5ZFIhyWol05h77u4FI/zHNJsLT0XOjnG65B
NVDUeKbHBEAsjT/icPBk9nC5nEcWhZRZzFp6FwQO6wFFXgpoOozZMKXB6NKfwvhF
iqxV3i8m6EtDryKGuWKVCXpaSsLfqSXt0cBOIhKw53k1yDalrl3p6geKEPAve2b1
uQsrFxY24gjMdXkBvT0JRfco/JcsD+Bsl+ZjpE7gqE6KSPJcj15IagdufsrJKw0t
qqJgCdvgeMVM6rUT5bJxgy4gBJHyu7XWmAWAWLKSOH4Y5WiQc3mPhZ4ujAU+iaS3
3gjsmKmmyN1tlYFP4CCbeb3A4VUhQWxXBhnsiz6D41AXM716D55p/mRbcL2ey+3T
wAszU5cZCwQBEgH3xF40T3L8g99yj6g+zBy3FTZRwIgBkVUUQ+2zhlyCpCFPJU1d
3P3qi10z63wAMYtoOVrPvNu8uSdoKdRwrtbKqaeNxirH7lpJrOvXDnlQzyWL49sW
gq7yjNUEHi0SZYT3yRUM5pYLXFB/+fX9lEsWRs5W/vOBYq8Ed1zDkmxWpRG9jXQc
tfYRUmGFHIOfZ8id6uZInVVJKwMoIQcuz2OdqntXCA5BG9X6VqYyd76s0SzN5wa8
nP7IE9q4ieP3DOGwyZrSgfmBkDUTkcg3GbrFOuIfNByiwXv75ol3yll8/bZUJH1C
H5oGNgSAcefj0IJ84LbtGrycrFw9HCKlsUW0y0SOcXOCRYqS/TxbLdfNYn+wDT3w
FXB2XLcxggECKZADxpJnxbxuW0yytMfkgbo1j1IUqsBJi/mCQt8ZmrhfT7V3BS/o
rN3BXZ8rWsPDRzYBYfi6Aci2J8UktZLEvam9sPPzs1Ftg6pIzU6fmWztQRpodwcQ
LGqekS9ThzgMtlvd4P31ATZ/V+1KvcgW5n1NckcQj9sD8Yl7w/ca8vnhZhAvsc0z
sNdap4Rtj2oZ1PwqecG7g26P/ILveNH+Jk7sPLMs9Evu2cjkvr2gllTn4UDS/3HD
DRUd5XywffvmbvLB2tz6weUBm2GApxnoUILE4maiI5gqmlJ0KKX5AMeK6c+MMPBQ
ePEak6vbugW0nMZv5a/regmiV3lpKS5iROj5Rv9TkltrWdG87PthtQGS0ur2Scy9
O8SDj1bKlsjY2dISq6phyVxtIIc/e663oE1ldJzEI7Usz2yVvgT4zIQBEj2pPKfJ
y5t69bypqugQ4dUCAM2qh1mW4Nwvn3VE5GY3oAiiD0z6SNZ/mtkhI/1uLMsaEMkp
AhQ6nxzEFz1TXWOsURMEPWsN9Kq7pA9CTDnDW3F2eYzPQZtvoiqRUEk8F9XTy5Nl
A2dezjRBSWFP+DG1zsXqLr/gHSX4277jDAjYuvejPusq5xeimhaT0vBawn3aVyy+
1oEGUSlzlYsfkoxzfzFBUikug0MROOR1wcWUWG1b0B+4msOQdO8gx6EfO6kna4Zf
d+VZgQw0kzj7FcEEZ2DSNklK3/sWIkKxYrG/Jc0G0RsIFBOqpV1lhi2JH0GkpZC0
n2K/aQvfuF6Z88ZDSPHpX6lqHKlKkSsscuwjwoQyljmggql0ROE6PYbkOjM7DNce
/yNaniP4RfsyCLgtO55MwKek/K0Er9xZJEJgTm3t0cbNRdmWl3oMz5sVaslDOU5R
wLHxWSCJQgKTfH8NPnW2RWDWdQURq9xu5v7n6u+qp3ZV7Y5a3hgAMrr8uT7Vid7+
FSqxMmniZi7r1vlwOzLW2PiR85khq2Djv5/iw+LepaRRplBpT1ESzyd4Q6RssVW0
kOI9HidVi3Fh4sgslNd5Xrw4r5wdftlj0TlFGNIa1coF3UZzxV3/shclCP/wAR3c
63pnM2JtGlmSsiPCM/XRMFgEoyC43OvZY9Ljnn14QRAnFG7/sBZA0GZj+iMm6IJ7
gpA9yJ8jIJZ0rQnq8uHj1vdSlELd2LTu1jpQjL3gp3xFsKGquHdLDWO2wKF0fyym
sYx/rRCwQWUfSu39U5H/EAeb4fsSoSBlBOCeKrQ1O0cWg86wFDoAbGqUi2EQLq9N
zm65VipD9IkqiXFlbT2Ifqx4nge+D/vLj0LsJxNSNr+Fq1e0jDXl+J8D1iQCd5zj
Q3KC66zVt+omg1kOCnekD2WIONfrF5iPzuik5wNC6XCiI7hmqQuko4KWJ4zbF3l/
rZ1LlDWW9mZtiyUSyFi0B6fitQ5phAMy3r8FsKc9RBo1USXWxAhZncieZcU09pom
yNWsOiFcX4fR053W/S3vV1WnMVgWHc7BqC0LAkYB20Zw8YCLDT+gk8XWfmp1fA1m
GmZF/EfidAorx9oxX8or6jtE8pwnXHN4yDBRvJ2YaXu+oZwIXyaUGCzwXgTDDbIb
LP+/hMSUNb7W5t/wFcxM5HEx3Qn2fdQXW9DBT0ClV3KVrJ6moyH4hp1vyhjXHKg4
6Se5Llnutd8mgfIKi9/+ytIcTsSwWvwmDHeHsa3ygxxUphQ9F8jHgl2S+A3FSWET
A07yZYbVGGzx7SyWhoum/3M7ZJUGcTZbQlAZQBjn7nKYeSrcZv1sb9Wal24JDemO
8MSsowgn+nNegbDXlovPosAtuJX0oxkcceRutlTlLjADCRwZ3Nc8thQNMzvmWSPV
szxVGO6XTI5IUoMp7cqbF5v3vJQQc5+6Fih2Afn2o+z4Qk6xBzMRQMZVJ9wgUw0/
+eYtUqV46vs8nUaydBmO4S6RixNQtgsT+qfWtvOM2QvHD5kNmgUdodnsD8MyCM4x
QRCD35kgJpAICEP26rKLOle5t+eWVRxE0yMDkg6+vo1UtQTliQ5xZeo+F+XOOJMC
hFQYx6jY7sSKZrezfaPu8pvZUvRF8QEOnBaAbP29ZXYCOfQT8/Bauh2REn023lxh
y1J5SnO1HXcH6ltsgEWMWszabMSRmh8dCsW2wrIxk+B785ez7etz3YDCLdMs3OjP
Gr0j+MbWC250F2aUuWlI94hrN8cuAZX0NY676X5Ij60EGKconGFRHhJ15oc7QI1X
FMGESrmwLZnBIBlNxwKyTF5wrVFqZ63ekiGeVjKxK9rsXxfXYQLElqsvmTp5m7Nv
aMSJO3tann1UzEnDf1gAE9nZo/q3+hLZeED845EHlu4FFBQkOopdZ6Or/I0CZ3cb
aAvLc3p2XP2tD9Ogbl7jXaM1uWDPmXHUdX6aOpmD+pHPZiBRdyWbNWQCQyeEtk9s
7hGRmCxYjuyljEKlueULggcoDTXn06sanX3p5LEfWG7sb/TxJxel6UDmNgiu/oOt
ByqygwM/D5Rrnfvyn3db976Go+h/ub+HNM84oy4XQPf5YQOFM2uvKdFnISG5hy5a
49A8/UKj0D5b3oOpQqq+3RONN2pGYe+kkzYJFg3vZlaFMMbIYKfidHajJJFtPGT9
r6ClNFS3uX5cW55CCOYpmKNU8rV5Uw70Sb8e+EnXpxLTF7eIL0pWciur8VZiarKt
dCUHFdfd/HVc+05vp/yT3AKX66wXEZ1mPRT2KqNkDsuiM0ofIQMn4lnFB2RmFPyc
JtL4DNLMfGSNstmiGBCYXUzPWIOTsVHFYUaxKCL3Qa1JJeFCYygYlQdwzoIbw0gI
LH8hQne/85FEf86nBeDTZqU9HWTgz3x7+SYGUZ/BfM/vpse33rqWwb6NTM8znl9v
g4cfHDE0SHa6B+OkIM2ejzl0nZ1RMVHtfDQTj408bRZ4lzQVsAz0RMS2BMckOrxs
bvB8cEIUN6sIG+sL+EKQfePnyIXK/ViEKlQfCb3kEBTsO7HLF5h0Nle0YWcEG3RZ
BGzEzIFatQTGjQMxNPyNupRmBw+X3+OZJUoCQSgDYZU1g8Ie0VJDKVNe2LNjITaT
XSf/Olk5jQ15kIka5oYwPVLXwmZiUlUQUg/9oKG/3Pd+lJ6TH/C1djGwoeIaeiYP
jBXZG3cfSig6MNXzJZQnSXDqQIsPrV1gGyBW8SKEQqjqQXshC/VzXDcuHq+1ROSC
/qJtsotTo5kEOt2R+UV3MpAthGElgB43vnRTwG7lFYV7vlYFD2iyyiGWKdln5hPD
Mu5b+lllawSXAqNuzZxbicqSJ3S1XQjRZtHJl7dyKf6sgQc74uJfN+jg66iWOqWp
x3Ly83Som0srAo15fW0tdliGhXm9dtWc7HP2vMtbJrgTsum5utI8qLQbXc/P3W8u
na37RQLURChQdaKPiJuAhYM4lLmgW8mXuCxM2uvmHkucqcqu7YXquTgDBkuNFar6
UOiC8SpyNTto7nEK5DWXGNRvnU2OHfcQLb7ZdKJzxeutGqwvZbznGDxry9p2OSJl
SVaWLjM7XURS3IIrHK1uEjzPgdFIgrlhXZnGcx3ZOQUaWoIqQ/SWBhrBFTIUxAfK
Mjw3SXlYDAE9fIPOa35BmGWRa8Zh7yM54YqsmRpF0qJKtVyLbiFKFW7uxWZWWWJ5
M6O+LVZwLn7knmHL8G2R5AdpSEf0ZRWIVuYGgy4+Pof8jNC5CEiW/W5sIEiqt++Z
IdM4VFlqAQFjlt1uoV5v348bxgw1AiYEYDYvr632Qy24TkPYRa9CL/vPdoVW49Mn
A1+sWegYFz0HxXzhQvYqqk/YmN0AYoQ6SqJUVZb+i/7dOn0ezbiCvoakARmf7Ulp
HsEyf6843hJWW9SGN5l56aNoK837LhdDpctKwm/HEGnyIrxVhXGbbTlFYRbrYmm5
qFv8x4NTFVPkmsmZgCjD7sbIJEH84hQq2boAREcIYn3i4Zqef2KrMO5BRftFoPi6
EmPkUOs1jxCFpFc6P7pojhjS8+OIDReRmhvvJ/I5pR8h3/NuJfmGmv/Yknl3HVqS
4zEsuz7tvmARRjY5ZQ2CyeYiNCvhts7/Qtz6nEFxs1SRccuoZqqf/qqk9riANBD0
+eFbkl9bSD8qKJmn7omI8RwcKvJ9iJg1rhWqW0pOMwyCjm/SV053Mm64woR0yaBg
ZUnraVYkXfOv49fIIay+oir/NsJnhaI8VVrbEZCY9fN0l/LFg0t3EJSBw1iCXAev
ZMjaOg9x63QLvuEbVs9lSyWz6wi0QjZNx7y8q8Y9ONI6D/Iw19UPY8wh3CcM85Nw
+TZLB5GG6OAWfAYqy0QS02EyrNFsPmIzGak3PhGS7aTgJnbeSoXCNQno7c3U/55E
l7kp5IqWrn2X76XgzHp82e+WJwgq0OQtt8enMmM3UnIY7vstd3Ct/9iUhNaPZDlt
kQNO55cGLVZsv9W8qNIEmUCprCemjn9UYyMZxXXBIbeQvNYrH75XknPZZMgs3CFb
huze+CcOGZN/sbXLTcaM5XEQDNNAsHG1obuJTqmvF7G7Ga9Jo8tLnakHjkGwMfbD
KAXPzemUXkPPZa5UqJuWFthE1sg9/L+VK9JgRQnC9eCMo9m/cOEQrAoxOSXoS6CO
xACGZZx4eEmEOtuaLhyTrK4HsF7TGEiD3S00pr9iRZw71946cTKWi3sOQfQV1LnM
5WTc2IQiACnm4P+xPVK7/PUYCu2uWQG3IRf1f6lOKpp/rVc1cNaMm/jleQ6cfclt
89cUTeuvmkl7PBnV4eYSvxmXMsX0UNH0DG7wFTtru5GU/enUkF9wKiWH24+MTEaW
MDP24HZZNllyjbU7cltEEkmLVih94LM/Awr8h5W02HT9AEJ7BF8r0RHemmeRcSvp
xMTZ0ys2Uze4aTVdkUMq9DODMgaMMQ96qGO0xDHHVHk=
`pragma protect end_protected
