��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z�V����u:0��,Lk�$�V�r�Z$ƞ6�xp���<3�k^n��ݞ��&G&"o1	��)2A>w�_L���)nJ�iT���˟�{\)�K���J�M�7�AR�u��h�[�BQ�T��
ܪ3U��+�g�h�	���g�D��Lŋ�^�`'�:T�8�n�����/�ϥ��#��'T��EM�RF��	� m�+<���u��F�tfU6�KO�~�=n��iхU+x��O��)$jVD3,%��h�t����P�X]�C����o�Ļm��9rw�"��k�U'�<����b��hv��!Ԇzt���
(���E.���=�N�"�DzhB��T��Y���-8�>9�A�&ԫ0����։����U�)1z�(�ħ�>�$�&U�xM����.���Gɔ�)�o���|�[�e�%�T*k��r]�V���b;4^G�J��\��}RL�9�z�cU\�BZ�Oh���k�e՗�2��?�l+�࣮�4^M ���Q�Xey���̉�3��/xo�o
͚�UPG�&�:�2O��k��=��seȦ��u���x������8		�>>�Y��w�U�Zw&w@6OtjO�'�@A6�f�P�F��U��İ�H@�:���|�g�rD��=�4g݉ܮ� +�S-��t�0C{�r���OL��0��bx����-X%%	3�B����du�`�hŨ4CS�|v]�q2I��F�]Q� ����Z���,ˇ>x>F�;�L�'E��]0d%&��{w$�24�7��&6>�j:�EU�]v��Px^E`�p1��1�$J����[���Ө�f1����?�~�2"���L3_I�"��X������|~�e�j�1L:~��:E��~�8W%n��I��q�x�#(B26,&�����SM������2%����d�l��1螦���ļh�|��V�:֐c`x⭧�)�߄�+�oe �� �c�����ա�:�k�Z��g�b�εrMgH<XVH?AHb�-�S�Q�[�B��q�v�$F6��� ��^��d���v��z~�x¡���R7(��o��w����N���x1D\�zЩWZ� �����nU��>���R߶*��H�!X��u ������ȕ�<F1� �62�����Wy��r�=�ϊQe%�?��e�ᰙ8.WS�mG�T�u՗���������h���g��.ش��??(gH�K�Ҟ��c�Y�t� m�ب�ެ��\�<��c�`�8c�:3j���WA*��U=�Q�A�y:C$�j(離tiT�1u)T'V�'��5AB�c����!J��l6J
=��U�Y�����|�-Tln~`u��l,7M�^�N�V���_�`D$_����B�#w�
fT�|��RS9@��[m=��"���`��U��H4!�7����vNǛs�����2��bW��>��b�16�)y��lJ�t��KP[��o�L���=����JArVw��6��v)j2���/glm`�	�B�t'&�Ϲ3]�����n���q'�v�ʱD���H2(p��Ź������Jk˿Wmy�@��3=����%���tc~r *�
�n�}��@W�^H�(T�K��D�k���8 ��,��x��э>n�^������m~�͓�R>w�l, �){{jBu�N����Ā�'h�K��K���)�@^s)b����Ƃӷ�oF�����ݬ�u���N4n�%v`Л��#���?O�z��6���o�[��,D�a
_�%���ѩ��V���-L�%8��M2Ҏ(�i1w�̴S�|���;�_0w\��y(�xʧ�I�ҋ���P�d1W�ft	*jZ]a����J{���8�u��z�n$`K�n����S��DA��&^�fCN������K\����̃�W�C9s�ը� �#����tO ���-'�A�LI)���!�!p�����9OF6�Lq]JQ�5��q�J�s�*�y��)�9	�P�x8�&�/�&������>���l���g�M�
�鋿���N�/�Y�q�%����*,��u��e�X젣��+5&$�LsH#���=��l<4"�
�����R\>�Yns]R=���Unc���V���ey`�u��KujQ++*FQ� j:��!ejr&������<���z0L�(K������Y��8�0���'�vʭ�z.�Q~Y��&�/~��=ۍW�;��G����ٌy�#�6��E]�Лm8�CLVd� j�Al���Æ�\SR�I��� ��>����5����EA�h��ܥʭ.5K���/�O�/|���h�co��keu�R�օg��&+����/i�U0�9�T���ٷ�;e����jTN���.@�%��$f�4���t��\^Dx��&�����Q�,��!��7����G�e�YP8���2