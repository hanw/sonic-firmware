��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���~v)5�'rs�,�s����kz���n(l�{]��h�+�dj!��A�����}.c��4׻�>B�ىg40gM6�݃�p�T�^1��Z�[�/�k�0lMNv\�o�Q��m�F�Y��Y�;י���1R��B����oXBHB> *'L��o�s$��1��[��v����݃�m�Wv��=?�Ϯ�|7j�u3�����͊Є�Ķ�RT??��_����$�\�Zg�`/��D%����8x���0�9�y<(�+	���y��F��$h�-���R�)�V�b��g��-����.�лʺI@��~z��|v��ɵ�tW<�S�JoxЌ�{�+���ɾ���
A�v�=��%��k���$��Z�{P&�e�uP��R���0���z�Ks:��L���.u��Z}mN{n��.+W�/%s�߫��`D由}څ;-<r�G{�3KL��p� u�- F��Q+�t��e��<�?W�$�Sq�a6�	`�K��w�{�����^��?|����+Ȳ�� d�h��5wñ��p�Z;2%�$�ʇy�1�J��8�-� 	�ɰ��Y�DZ����ٵ]_*pKz�%��Hc}�[���כ	�]�\T�QSI+A1b��rW��Nw�E#���("�y>%
0���q��j�ӿ[|�hV�!Ea�\���Qk
��♿tq��!̆��~d��A�E�y8��om<�T wy⍺R�[U���yW}>;-*�����Fb�N�v�;9���>?�	Y	b���v%-���+7k$�����~���X�)�r�J�6���T9����b��^�:-w@0d9Y�b�f���� _ �7�oӂ�R8/OsǙD`̆��f�L-�:�!a��K�cɤ����P��n���Ѯ���熥ml�	��I� G@���Z�Һ�����j<�.4WR_]d��A���>C���~�n���VW�S���Vs]r�"F��[�Jo�����e�w���f%c�2"�D���R�M�f����@���5TY0J["��y�eV/3�����4]<���
�a�L����^�҉`������|�C��A��K��xQ8��2�ϫ�6�+�ed�M߁*����ӘGOIȿ2 p�Y.��FBK}?x��ID���f�M��Z�+]$��bG9�Zga7�.�GКP�]]�"��_@�Kk��!w��9�`ޣck2���dg4T�dOF0��R�&�E���w���d.T�Q�>���l���W�Ъ���@��i����nO~eĈ�-�}o���,_/��e���?��9'��^>,�Ʉ��������TԐ�`����[�"Z���l�R�� �[���:1Ede%�!��6\�F��2�+Y�T��}�d����1�l��Fxm�+{��^�]�Uq΍ ��O������j$����af�B^�M�E�ӭ/�a���"���q�ݨgUj���Ee�o�&D�M��m����K�V�!��%m�jG��6�������Y�Y)�/t<Z�[��Y�����bND89�#2ӻ>��(�|�d9 r���V��:�{�� �i��{iBHR		,�e��H&�p�'M�!g�9剹K��Z��|P��RN��.�͠�T�r���Ϣw�x��^�țW$9f ��.b�=��Ӡ���j�p�a�طl�]�O�1�dqcz�'�;�G����o	ۚ
�h�$�"��\�$V|��	0���J�C�R�t�n�)VI�����^�C��7����n�q闽.�F�g6�@��.x�1�{��hs�<�Bݰ�Q.�h���B�ʑ�hi��z��k}D�������i-uS"d؆�����i^���RgU
8F��7&q�J�L�����\]���l��{��bA;�5(	�hPk�#�ۼ�;pF���/� �#2G�L񑖮�^��$p���.���K�$֎��������r��ז��i�����7 ��w<KO��r/�ųz��B���tP�
�6�ۑS��ZՔ�H�k]lZ��o'�l�(�kH��~�� 'Ef*%�d����o��N��p%nw\�;���G0�C�"�`��
O]�\Ƽz�%QLP��(f��C�01IQ�y��̩�����MT�l�D�J�i��e]�!Q�����Guߏ��Je�;�{�z�i׷���ך R�� ������6o]���*?z}��:�fE�w��UK3���p7C���y�������o�b�T�f�vtI��t�E�QU�c=>þd����E4� K�����@�J7Ē������r{�$�����.���V�	P�Tv��?��6T�+�K+�p�VPw�^~稔fҫ��P��,�Dl-ϯ�< ��N'-qo�$3�������b�?�S1��7��T>�_�(6�Xy���J��Y[���c���I1(=��@aq�8p�Z��޸�>^#��8�$�����ĚbJu_h���%��0o^�ż��::]ͧ}��3{�t�iIimWo�P��|�����Dϝ��%�ڲ���y��x��p��/&��Z�B�Y���$�20��Ɗc�;
���|�������baQ*�	�=�Is-&ܧCw��b�7oK6F��[P|�,��9��E�Q���HVn�zq��d{�صђ��K"�;)�F���2	6����n�=��B�z��h����.Y�}�S;�CS�i����cO5Gm+�v����|Н��J�Z�U�v7qQdtW�\��?ŻY�L�'p�(Q��B/b�D����~�I�Ë�G�U�?���@L�/���˛��
�DD4�Qb<RC�.�}��:}%N4ބ�?��&ޜ��蘝��:��X�: )n��1a���ji[K����)VV�V>��k,~�bo�<p�ռd9􋗺�mn>Z���+�B�T1����`" w��8�)�k�n7���EE���MR�:F�t0��B�'�=wE1`0�%,������ͭ�&�-�r2d���(R��'? 4��� �bt�Êp��+�׀�K��8�k�u|\��w��#�4��ٕx����z��n4|yk�1fC��Nv�]�K��K'R��͋�5]M��Y&i<������r���@4eQ\�UC��_r���#˩�{&̃"�oV	*�mb�K�
*���Km81��a�Q��i7.NlG,f9P�����C0&��Ms���������b8��0�@��bc��~�̯+Շ� KZAw#��(����~�����%־��f��������2�ԋpOQZv��c�ُ/�8�p��H;��R�v���c��n8��h>G��:��2X�	G9��er�;�?���8�&t��s�wru~�����'D?Y��iG���s�%�rбא?YxW�	��/�O؄����z�`������U�bN>*�P�Ȫ�
�Kg�.�^6\=]8��<T�D���ys2�9��b���o�
=�KEݦw�p]���{Y �C�q K�Jf��C��i��Ǫ�e����[(J���@m�~�4��U͊���1 ���R�|mŪf�ر�v.��Tb�ݡ��Z=��#��{������m۱ף`La0�!��U�^eQ�(0h	FLދ�I&n���9\���%��jL%�i���A�P��%�g�\�;�k��/(1K�B�cdq�z�I��`�a,���/r�̏�%2���ӑ+a�/�ydܵޫ���ij� G��^�?^t�9I��nX@ ��oN�`cS�cm�TH@n3N:aaZG�Aӽ��Ş�˪���D����BEAE�h�y�Jm��A�w�|Q<� �����uXk*]5����b����4�#�g..�'�#9:�!mu��98����b
���'�7�|�豹�������$��a�Y�d�ՓC̬��A������pin7'9�������qT���[(�#I�:ћ��VA-�,8�HP��F�����kb����#[��>��P�[	+�[Q
���W�R�}~� LE�Ď����;i��K%���1�@kո�X���>P���I"oa]I	���n;�\����&]�W��0A�/MkSa*��].��o�j":�;	��VYb�j���oe����6��X�<��9ǿ�"�آ��ct�q�uP;V���<nY~�f(P
gh!��U�6�ɀ67�C���P �\�'#O��"����G���yT�$V�^2.��� �RYfH&H�oV6�������^����2)W�
�]r6'��\BK�ɛl����_���9ϱ�t�6d�{W�`��8�����w9�Ʀc�X2e�3rJ*m\VU\c4�!��c3�n��މ���}F��Wh-��h�+����X�E�9'2�Ճ��=�u��wGn�b��ʐC�k���:�-	Tj F�UR�(��by�e,���Z3{[�X�Ɨ/͵d���L_�: �&�����s��x(جnsY���#�(�Hz��-�`�������*���̳��c��PoMX�=tg�.�\Ցi�[�4���{�Ν��	8�0�X��d��!�9�Ǜ�����+g��c����&�@�oO0H�A�/�>�`��%�*U���*2듾�3��	�[�d���A7�צ�:a��j��sb�6^*ae=�ԣC%�9�j�İϭHG0���(c�x����
mw.v��E���z�c��ߍ��#�yٖgb�#���� }�E
����!i�5�lhnm<�x�2Q�_�r�۷��t+��WrP&�q�����0x��v�{<�� j��V��9:,DP� ]�d��j	��j-��KT"b�>�U|8������9�:~s/q(/5L�*��eM��-ݘ�)��� �G���K�2�3����ŉ�����$(�&[�����&��d}8��/�97$GA�Y���Q巯̝����&�p:͉]��z�H���h	��Sp
�:�+շ�� SZ��S��2`q��m�Χy<s���+@[�Z��Q�쪧x>ÊO����a������L�v�O��ȱ��1�S�)��˔�Kǻ#52P?��G�n��m��s1/��s�����hWW�!�a��]w�Y}�2+�a�b�ʓ"�a|T���ӽ�������2A�L���7�Q2��'��52?~��zCѷ�  ��?x�[	"%��$Қm1���8[��y���ɢ���^�����[<H'��e�C����j��VX�¯"(�X�K�T�lm�p�f��R��b�N�b���"��g@�:�k�HSa���{�Ϡ[�Q�����x�B��Q�"BGfJ�A~KԌ	#D��--kR�5;[�I�p�C#U����������� ����\��I_|����6oY64>v>�%�\|�^�d���%W����W��]
�6ޒ$�	c�A&�}L=(��{��ׅ0n�{� *������m_���Ѫ��̡�]#GX�)�|Ɲ�?��5���S�׺��}�᠃l+ͤ��&��kV0�r��x�#������7�T �^y�p+�V����Y$�tb�.U���.1G1��؄�G� � ���
��[�|+z�A�k���wE��~^�o�9P�Vx��K36!u�{�J3A'��辑b������������#����3
+���U�����j%9�=���F2����A�3��'�dX)�
��M
�p��5��tN}��ɘ\�)�&p:�e0��ߔz��@��yfD~�˫D��\��̳�u�HVHx.O�y��v�UG]>�$-_K�U}�2�oM���C��z�u����oW�D�M�5������8�Z��"�J2|O����H���RA+#�_�I6r㠬lq¼�����Sa�e�8�T�R,����g��}�����®ت�v�F#��,X�Ì?U���j��ׯ�P;�v�ϲMP��Li�e�hA-��M�;C^
.)����l��R鹭#ߏ�߮�:9�YG��Q��p�V)SP�Aʈ�r-�FB�#�`���ՙ%�y2�<~�s"2��W����LSH'��xǗS�i�p9E�/��y�Fͣ ;�����x1�0-;�����gIFBnR�wd��	��	��wu�ϵ�A��^�/�	���n�MNത��۲<�����!"�l��F(I'�Z������Z�P]΅�o�)]y�_�R����̡�8fdn��V� �_0=�X�ͭ�ۦ �gڀ���q��O�^��T�
��9��"KY��"���~l0�tp�S�+�E!�埫9����!R��0�*�rw�'�Ϊ�1e�����E��M!�F��N��T�V'�A��t���Uq��,'��j�ӆ�����j�1לH̯j��ϕ�|A�)���~�P�Q�����z��oN�X���nQ�3�4���׭��%�ȣ�CP����̝X.r���z9��}���;>$�dI��»� �$`���� �Q�ױ�Q<gJ���\���R��j�r�b�gw6<[��N���״�������3XJl>������ے���]��[I��_lf$B6\ �UE�P)�X�(��5?pb�`�cL��ico�Kw���|P��E���.h�-�1Y�
1���O��G	)5�ut� +�2����j7�r�B��%�P�Q������NAw���=8��V�h��WH�����B�~w��Y�P�D�|�t�T�%-�$�{5s�,9��xdGWh	�eqH"��u
���G�pVP��V����&�1�v[�eS;9��%�&�Y����qm���Y�`�!��ۓ�-�]td�=!�K��γ��w���u��K� u񸵬��wG#��[�^']X��6Pw�Kλ�kN%�~�)Q��?4�:���)�OX���q�px��홂y�O\5'��s�
�3�^i٩��#"/�XG�!`���`A����jn�ɺ����)����,��:��:���1��_`�9/E
���z�X�ަ-�Z�J��v��e��Ϝ�����2��Nn]�ڕ����%_�Pr�6���U�x>Qb�����O��<�>�us)$Q���{e�K�:��#�n:VUv�
v�ǩ� ��$��Q�(;�;�l�<��L��].1.;��+5`�3y�>���H������S�������W�����lʊwM���e�ʘ��xpq:�||Hi8aAa��K�$��Ob�Q�[�.)�o�ع�{w��06���a^��yk^:>e:pHjK�%�����Ta��&�
M%��z-ى�T��@`�Y����$S�p�S���R^���:������B�߻�<�D��**V�������rRrRI��*<�mO6��>o�ψU��l�^���j)E�)I1,F	�񟚁(�!J��TM��hf��k�q�o������3B�g ��Ky-�{T�Ż��]�A�F��:њ.N�d/!�d�������&�gT���B.��Ӹ��"nL��A$0�8Q;���,������L�K�I����Y�[���̙�����B��㣝�+$;��M*�����T���R* ���:���I���'.����
��n4n�x��2���_�� ��C�{$_��]̨@�Q�(��L���]1{��y�燸Y��Oc��G�,hXq8�c�X��A��7U	 �s�JǸ�D���ٰW�C��p	Cq��s�1����2k�'h��ݰR�Q\R;B��9h�"_� �P�<N1���(�^��6ݜ��d��
\LG��6Ab���qZ�ś1gy���7��lO�H��1"B����e����d��Ⱦ������am��Z;�M�j,�!&x�E�9*ozL��z$���LJ#�Uz��-��M��c.�`������3H}�jw}m�a�]yPmXPʝ[�øZ5����N��M�(|�.��~����퟽�~��	��t��|jD�\
Q?��J��ׁh�weW�皠Yd��嵵�)y?�ێ�����*���0 ���=�Vk�'��Y�����RV-��3 ��k�v�Lb	��bQ�M�H�n��#,��o�e�?�q4�T�����A�Q��٧����7w)1Kn���fƪ���:{�x����"`Q��$�^Wjm������4n��E����d�J�`a�8�s���+{�³D�E;٦;��-z���[�^�P9QN:�)�5�01�ӑ���1�/�ڟ��Ra=ǹ��F!��|b��F7m��B�\Z�h��Q���l$���\4��<=Jݴ|�J�˿.N�m#�w`A1²|�8Q�!��L����{��81����a��G%�4�\��\��)���?�KE�Ԡ&�O�u�pt�0���� h^D�eӂ��1��w�M7������z0[��Jbj5ˀ���,�!Q/�d-+���2��Ԟ%]KS\�ͣ�jc)�Nu�j���#�2�p��G��.�+YJ
���8������V���T��2/�K�q��H'�n�FpU�.���Kn��n�޹�����"�#�v��k��o����)���A諳X�֙�I��̳h|���j�A���-yU�&��2@����c4��Ť�/