module top();
    sonic_rp_ep_sim_tb tb();
    test_program pgm();
endmodule
