// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
beWzV0qayW+N0p7NVbyuu0LPSwpAUVs6xzlpGpC5U/qp2TXjnyZw8Z6k7D7C/dAr
+rma5FBdn5Tm4AGeCS6MbpGgLbEqItRtRwQ5Jqm/cAFNFfoNX/D0hqYjJztEx7Qf
lrpAORzpB/B0IiXpMjLMEwIuTzs/kgGIiAvqH5o7z20=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
+vpJJo1K1UhI5Y5nhy4ixAWZxltfh/Mtp2G9y4PmmiyDHqq9j+WfKrmLnGkOwgUL
iZbgtYwEMwRMcuzRuexg+49iEBBWG4buWnvk3tRxpU325vVVzvXi6ZMobJXg+Z/W
0DKmdVxUoV2x/uAU4rk8f8XvfxqWm/6ctC7oZVTrb0ISEVkJ7xatA2ylM3jL8+Ij
ud9Z+GCKiP6A9oTPsQk92Ar5gnF162MXBkKD35Z+JSYLSVEAL17pdLyB+MucZDTP
bn//WGz686ihlQ/rzOwAfaB4utCBz9qNWG3RSSYgMxkvjmGx7qbV6JHnxqThAWFf
s1410fh//kAOP6wztavOsbPKcZ0ZQOz9+9COAPf0H0YGUmGATNMKuHMcf4d0AuE3
8oPjumdzCaO8Zp5tqvWeTul0NG+DceOL+mLYry1K4N1uK2u9bzq5N9/dOVV/uM4Z
qJxRgbiQv2lngMfENmXw5PuHYLfpwS5bXTjIYY99WjWgoOrYWkPfRheFAZG+XGzq
VBMSfUWL4frjPHs99KiYcocMwV+DrRfpxWVzTwIxIUia2ZP5OTG35R34W93FTz0f
nn3q+UcRFE6d8UkstqMixgDx4NdUYhWcym91aBwifTX5pPDqbKklEC+PC3bfaMVJ
czFRimSXUbS2cYk8Z/JuCjUufo8HGk58XNyZM5DhHaA+kZxgQn3NVqdMKdkbu5HD
YtIfvQdfmHAkrErXmHsUufnpYUPFBUHzPRt/S/VUKGpJvLd8awuao8t6Ys1sE7i0
WYGIsslhsAYqdjrdfM4Zt5RPV5VdbHP3R3WCqZjJL1pUW/RaQ0ymNvOB6XlCOsN7
Yush4F2Zptg6ElO8LOEGqRCzfVpqpHnAxbV3h1lHGLXGP5OXICHVXkZylOEyLWVf
atAw2jbzd5vjTvKMaNZy9EH4LpBv3VlnhMZT2QUtKKQU7llYPeVy0uJgQnskx6HH
Hsf5CYCEYS+7G0NpuBWE2Wz0N+6Wd0fKQFzXBo+mN58N2keJ7/Es5vkSO50H02Tb
wcCaLeQe6107K8oIaIEXJAN0MGJSnM3EuzzdGC5PP5pHmOp/cU9aPib2UzYqDMFm
3F2P8dq78nuf7+CCudOeevxJThzHlAIP2KudfuqXDGXdeD5GG4QYTbdw/yNVDqSE
q3OjZHA/pW8lqIPPHJzfCvL163UTQuFO59cBij2rnVOaS6UEhk2XHBVQUw5oWvdW
XmOfa8de0aBwP9oVFYySrpBXO225j6uF8gzfpxOWL76UzSxwi51PLAnyNkpw3jyo
izfYW0/QEkV6h3HuyMM8R2zyAQOexfFk/9hjQ4PsmHxMVTj+kwiaPE8rgeR3VYbE
7pvBPweV8oOndttDgVDExfO4jnHC8c6IZa+gfhue9IJ1wqj5pyJsON4staml98xf
aRt4PsqqbVQipjwh+bUh+abgFyRWOdIA2VG0qy66VV09iNtMN7nVbPIM1W3tftZE
uQZhyw15XRuP0RGYAGZk5PBH6c5bNSyQkdMO/wXAgT9dZILsSo5y9SHDf0ixUxzP
S2lWyGjLbEemhSBIBm0YflamWC2+Cg6DWyLmKJi9EUnC7rdsvSA9CiocsBLGHA2c
vMvvJyBBtV0hhir5WlTHx2VD6YQnFkCknZ+OoruIVtNTwO89fjMlO4+hxU94FsF7
fzKx3DSA3jyIB9uI00WpHxJ/7+cXC24gEIYXkiJ8/grCc28Y+60P75gvNLm4PNaA
NbExvcGCOfPA5aF3ORCB7E3gG9ca6nvSLkiwJCtF/dLVS4Yv0UEhB9x3VzOl8Xi5
vm/8bVGufFGmER91c74lSWf71iIWjxJhWYxHHP6VlmD5ZJA5ZpfELpt6v3n/fMf0
SGOYDZI7Vud+fXcgi5QGrUZpWGqpse3GX1+sws8k9/SW3DWT8031qXeOutH1u2OF
8QcZcsgebgOmczhdeDlpAHa4+7F8tolLYsPmewzcgrURTUa9UXmogECFdcik7921
FAi/iPt0xHGl/YZ8N4lPkyA1TGEl/NiS5r/Zj7jb5FdvAfX5QjM9kBfhXuEhU/Wc
iWi4cz1D+ngJM47iRYe0+mteXYaON8S/+EsXoHHrHWbyIknPKA3PwFTxIZK8b2Sf
h2L5PA6bqm6NThaksPEKLj7YA5FXH6DaufwFT1bx0s1puUWKeTkigVL5gmfGg2yo
8oEdrjrgWod21Eq3e9Kff64v+zbPgzNmaJgSHjsWbOfly7tbZuRt/J0+wJpw2yx1
eXBsZEyfCzkrKCe0C4JZ3rxz0gWozZdhwyWhMky7B9wxxyqV3TRyU8qtsKz3Vx9S
rOYA4fsea9PG5A1iH0fn9pTeDp3AP4Xu/WONaWUyrb3nB5P+gsLb+tGfR/D52nHC
5BPNmAYMkiTaFl9T4/W3iy4hKujIsleogkslZh170b49d6/vRG75j5e3N55eMQ6S
JZOEcKgprNfOAueVUgJ4J2pygb+18Z9WKiupOzPW0BVgXgNTMkgIM0kK31QDGT0l
Tx/pHw2Pwck66milzg+Jjpx4zj6oIUB0+/RlfPohHAGpxhnNBe7tbMlKYB/j13z8
RGWVHKjQGh3nUaEpwYsiQyDNfUT3wfWrjy9qRO7Hz9v3MniYHlfYZZRpIfUWwU4o
OPLyVEyT/57IqxVz5c4wDAsyuKmD+S4TPc2RbbAUe34D4o7LejowhLQoQNgco9Hd
7tDty23VAzmF7DU1XcEhVyETsJalE1YmuRPWeUSOtIhIfymAUiY0I7tMFrB0Mpap
RbprJgsXlm87zdmJH9YITBRSaecG2dZmscQ6675fwDLt9GSVH/AxiLXYyve1je4x
G2Bfip8O29x+q+4PqyU0t+ZUHji0XX/s8fmNr5hSi/q9SLwbvXNRMOTw64uO1uzB
Zeu7vVayP9SbHGuQ/E9kLru+fNu889s0uyZgU217IjraU8E4K2OxTEHnK3UiFdH3
yFKeyZcqkqy71EbObX1iP2LxUbPkyB/XVV66tav/xyGo4bKurERfwX45LRYnhDHs
PJFXeZRz4bH6y4H8c+7bEaTVjDLY0YdT0yWWou0WlZUL++gmfeSI2fF4hdH5k6CH
lWaLUMu83HfQxTJpw3deIMwomTGlsy4/ngMUacI86+MxCd46ZjM6z+r8xzIEdIID
srCgEnDrKBSIFAcp6I+KUrF4pP+gZ1XGdeePqhNNgpemCRF3RhGNhScD0ZbBLQpI
xQBBPmjWBCQwju+tfC+VT1dJFQ7+c4BlwL+ZcuTq2ZA7+HGvNS2mIwJ1chN7Gkvq
jUOUpiwsDyulK9srO/6qcg30JR6JVMiH/kYtqNWNcQoUlpOw+0ZcYunsn8YN4ngi
rU6ZxSv3IGjd/mc/4RLMx396WfH0CIhDEdoqEdpCjAmKMGU9vSrHs4Dao4UahZPw
+5yFoN89mhKRcQ2Ly9KCl3vikzovTDafsYl9+9cyjFmEWpuIYkOM5sObzT/xISou
GNk1nsnKDUnTn/7jHnTxTxnUgz7KBUK+ijvK6gpC9KWNds383dHsZtLdk8nf5glD
hOOai9GcOYDNk9MNMddrLDk2l9n75k+mSoUklEgainnz7ANB5BvXHpJVbucXbqCP
c5FLrpE3CkzR4iUrT+lUBn9ry2s0R/26Bn6RjmAMTz8NJmIEjRKG8nzQDQqtwpjQ
oXKN3U7MKRBO/pUiAKmIIAYbsvvliR0MvPfT7e35DA7Wq7LfW/Rn0AvrsEwPl4cn
xsCFScVlnIdpxv+bloCxCmsZ3WIlJx4obnAM20KNtaP+05KtYpSusO7o0K/MEuGK
kcraJODOgIm3TBFgI1vqvdRMaMAdATgECj64DMXPh/tKzZAwL2E3o0OHGa9cRNlt
KedbUjDImvfnIu825A/AIx9nV4BQ2nOPtZPeEqlaJtgx/x/Ieoe+ksygsNA77Sng
GGer+5wQqrQosmRndC+7p1zSKVZGbUKfSWC5gMpvyyzrYl43vTLiOWkcDil5/YJk
lVdP5pWeTsCp7X1q0inuwUdSVh6/0x0+6r36UW+OvQwxELqBAfmWdnOV8MHB837x
LP26Xx1RegBGvZdhmaaYmHloY7MIn/7fVWcRG+PM9/2MkvUp1S5ws5NaQV5B9Cqh
jv/hjPt9oZF2hDmKUz1uP6Rc91Tt0IHOIZxVOXVoztuHdVm212qV/boLYVbgRe+U
U2395g/Wrccm9UP23+/MxglUuwgC8iJxBXdWiFD4P8aiXJdq5yI1EIbylGe3kQah
U7oXyholfoL3FxoZ06nbd++sKjfzDcEunPXP+1vi+sqNirX5oq1+J+Tk9LjCfygi
kVZ1kLWInH3L6oTyxGJQT3Mi4HDhDubmPvb1pjvwvmfM+54OapLwp+p5MHLJt/XY
o8FF6T1rCn4Y9ffVezVot/6BrclPD/SVenrZvp2jw4lRWIHd+iEDnPYt1WNbmyuj
Bfqs6FAdpD7JExYuzMf6bTLjMTkO46XJzZBTxNmse8PHpSFOC7XOL55wW6ekd4KU
GivFdKqg1EfStZ4iT1KK+VvMOUDB8Ac3M95rZy5VuC4DWbvnMa2Q6Gorqd6C7QmX
fa6yz5HnaRB3aKPI2ZT8aK9e1YbYjV67Hq0JE1lOske/IJCTtOBMJb1NHj1LyS/H
ksPx21YERrAZfafm7FDAGAs7HW2zaREB4HXymJ2j7AOqYPVE3SlegmAq5X0HBeQ4
uO9LtZCdFVhBxUHrxalBRUD3k5g5vr/OsnZEytLoe+4r+xe/xWQqQRZ8YEaQO7rM
LK4YOTuOxZZjy0PS1J2T2aazGyqtRsU2WohEEzKyskLyP8TrVYpAlEsn99NQlP0K
W4rqzqPDLAfCX7iR5eg7qJizYUREYGJz39RC/R0l271YLVI8MVxlytEBWtC/g11s
NIW4F8NGI9YukZah+01AIU7UL4PTVK+6doy3kBkMAow/XY1Yfp5oFdKNHEjukdkP
IlHhrNQvSbgW0sxpYSfJWO4BmT4hUPdaUmeSM0egIX7ANM7ZjcamQdUfikw9HT7i
Eh/grIEY7ylpXvyBdQ02GElSneiMU0LoesEyedeXtUpHjumVZ7IR7AsvBo0eR3lx
EbPcqMiZefEmTQ5/HfJJEb+IxPgzRxGVIa3wijpUmHYLXiqaDEB1cAIJ2vsjG1BA
4IadyabkJEc8N7hzCHyBvUG8zGp7fgW2q+yaHLi55El6LwM9DwCgshIZPHSEL4Wu
oLY3lJ6SjPKGJht0rL/96pYFkqEN6cu++sNg1XehtdAPjnEY4OX3I8w9eO8liYkB
amerFA+Oep7H9tWA0X/Z9jGlo02rG5r9f4VlmfQEJ7sqDnz4QRAyGIDjkbdnRJ7o
M7aAoeubWrbj9AuIQPEyYQRfwIvRvVuLU7NPO8pCxTQIP1QG4gd+6T25OC0AsR0X
htFPIiXitSHWaqTwImu0QkTpxsFawO+j0yxjEQrC1ewOloDOU7TQfCIfGoMG8OW2
LQW/TaiENDwOZ/fsPhTwnSxFzBo2wlHZeVmcROx+bPlIgB9XdLsTLFyPPqjH9OZx
BG2X26TAwG1Gmfgoi6YngYN+DEmNPYEEMl8csBuT+dVOjA71sWgJGrq1IMbcdcQ4
w6SquZ+T+wGIF/wlIW7US74pjvIvZFXnUoHJtQjhvFVkHUUkUbhfOEl9v8mPWyNK
5i9Y7g6ISsTmpsJK6M/YUq2zxJL+fBpKn86CpB1cQGlvIMYxkCBu8TT2rLOrdmtA
DrzXZXejZ0b8BwM3MWW17qZh0R5xCJozJUQ7cbQtJbz/rb8ulpG7Y0BJ8mi0AZa7
RqXHYg7Ev+cPE+COImVIc/JtZGxiUJDYXp6S1C38q2ozg5/xQr0y6ag3TYVTcrdf
6ZAFukR68F7nt3gMA89SENt+HEJa8f04d1+j8vyNbE63V/c+lxlvjM1+WUZYL0Pd
9PpVWUkqTin9BSvx0tnEvfTLrEjXRM4B7RR2ijsHEYgYU0U3N61wEtp0wqQy3FX5
gpE/rKZyDGp6bvHtrRFx8R0NRUqiAO4Akx2x8zZTHiV870sbWq4G//t1EQay+zE7
mh3P1jyTcX1+LiWg+wkOhqNgjBjN5AXphIQstQY/8k7mgy44Ou2d0hHWuvXIDuLX
KlLOwgiULyRY59ok2K2Mq/d2joL6B/7bCOk71S+6E8yE5ZBSjF3ETAoXyV/AKj+H
MpUGjT6gShQS9XUQRh4JkYjTRX/TAxXG6gL25IyahPrC1xvcnN78O5aeVMjhpqCh
Dimg7n3mb+vzgcdMawKZmsmz9oisKvrT/rxKBRy1E6u9fFK6xrkOvH+779hqQHJf
s9t1COfWmPdnAl4d+nM/FD0ot4w9Mw8SsugRN2F2WEpZ3GdOFAsdX5eu7ysA6JUJ
ftaCf5r3BEytQ75Mo/REQdOlcDAcvZo1bcESeq2rmsDyVz7jafbbIHpyJ3MFimYE
eFnyUkLbabL6w3JRDGycze2ZlZvpRe52KP2546n1ZoNxeZVegmXjt9AFB7JDZbK2
BRQTzEKkYHQYbc2QJBc7qlWorpekXg1VWlP3JSc4ikB0gH3nAmwnzUo46SiOHiGm
KLe924uF2BL0K9a+BQKYX7gCrwapq4WdkJb+pP+X9tXeQjd7HE3a9MdZT+fNQLiB
piSUb0n+7a6rp84FpGxY33lyc7TfAttmcrDGIj1wYWRJLv3ePDN00PbncBOEZe9Q
OBSVFxxer+cm5jg3lotw5HwHZABK0yj5WKGmRqpI9bVwf+S6OgJdIKmYqEKWsGeR
8aUy2rfnceUfrqz5eufdWRmb81DAXKxw4o7OK6g6xWeb3MgU/0L/1VIoqTKQMc98
3LFpPqHo7bUv9CEU2wjrd3gnOR+u7eT/Pb2q9MXxO/PuuWObPU4XmEvTZ5J41V5U
6XHqZJR393SwAGIL498VOctr/faPECz1DEnIad8JXCM3LGZDgtmyN+mIpuJcwyvC
Pe9ng4jAvdxEm51RgoLYri5mT24pafB80q53vu2Bn1SBO+nVlZH1wHCnNCLXqa3i
1/sR58Be4vefPz4j83QZNPkoUaiqSXNV8IySo/8g72+AV5uVsYmHmG52GaE7z6Gz
cNGAWD+Z2hmOYRBNS93F1SHR0NdDBCsD4TVb21Hza8WPW6UmR9QHOx5xoBuJp+2N
mtgPe1efJDCNSbWmJG+RxDfkYRj3Zyh2TDtK4wQe3qU8IockirDlUTBfZ/sT82CU
oZzTtNhBPaWzgYtjV3Vtaw9/S/lgxu6TQGm8cj0E8mYy2mC5WkIaOfkrsKbmucyQ
o2cbjOovSixv+vtvyz44HD0H82MeiZzpOF75EMODrXYllu+Kb7dZOkJQ0npJzAh6
ajQcCF4AthHeF2pmtahaB0AriYn8edX6LO3q2zNfs1Cv/DKx7KCTtUqgVq4sSDs8
9Rm6YpCQHUV+JPC8e2ZRGCTq34eICdkgb6YXy5QKrOhrCKNYGk1l7wTFDBwh6zFz
ZN1M9cczGAV4M9bZII6ybxazpdJNga2NattdurIGsjYAMXEI1hjb2GWkhYSSnik6
4gTpCjmVJGYTc+MQZDS/J1Jm2FTzP0utr580qYESeRWLkm812HqgAINugWRFqM9S
5JodkeGL/LK6t8VTh/3mWaGFT7cwCoGTxtK4KuO2bC4HtW101u9LePA3vu6gvtZq
8ABnjJchoddpkwkP9drlHC7o2i0lyT+ejLd00UwklL1VbQSWvt3TxW28X3mPdUdT
9ME5HHSWGxAdHSU/s24KXmUk8G4iXf2GMXRjA9G3Cvxy3sJZ30fnYLuw1qqSXpDy
6I7yZUtQsNskcA16Uv3nJT9LHCKDyF/jLH2L5ugwktwzWFEAfoefZhKeOsmQsQGf
o7/weLJ4CGlYzHox3g0MuiUDMxVEApkoBnrKVkgQIB/NnRDvBFDJvgTqTR1dZjvJ
DopLcGwl/L0X1d0ZRihrUwU3q3cr2I2ruvOAyNY6dsj3yu5u+d9ZVn1P4r0t2RN5
Kr++J+vFkn/KcOU1vm5h3WjK6jTlp6yi0BygC/LsbTsopbEjwBSjkyXEwIdLmbI3
Ddtvlpf11Yet/xn++PyC+WTvm4ftq4+jf9Rbx0uRzDe1K2bX7EY2qDDloFoBq5vV
yFCmjeFVlUN5N/5OgHJwVVIPgrZUbxrusxni4P8U+1kI1jtef2HqkjNvtbi8vxKf
m5hGdzi6Zzqo1nNx1JL2g5xrT//lyZuEzVh8AGv01+FgBbs7D07GYWwh9OxD8S0n
fYeBh+evTlw/0onDURlGu/QkQm4QjcSBpMUnd6p6Dr/PWEOCU4AaKznjXVCY3EyH
WrnphxCdyunByVqUt47j7oSK/wUX0J3jin3CBDOpFLg6UFHFNChsYBC/IMvnd7cG
/s4VEOkCKFec263cKmIwE6KO/7gMuhTWT/taKcBRuv+rL54cAOH6L9wez8m1wlCy
6PIXb7+PMO9d7R9BDdB1d6BdIiPr+fhu8La9Z1Nds2zxAANIFiQTZbU3tsvEQ6eq
FauwMR88K7Bhdn6i2K2mQVtnub/d9a126/M6PyNyb4LlVqbqDtZaQrtfTI71x/hL
WZngvw6c9UHBwwM5MvHDl65HVB/s0eBtbckokcpxoHDWtLc0BtH1eREd9toGfaWu
Tk7pYjrOKJifCNP7hv9qZ3Naai3XmSNCe8wk0rL7i4LSW7rE1IjpkthtAZv2FO5e
reptoyF6wh1P6kWKj4FsQo6FOS3grOgjWOdVNIsjwLB6UStSbqaOzWAJZCiuYuOp
0mYWX4f1yXBugDdBHeNHg20vfLQoSNUq2DnxvqhsgR6HwxjiAZccaH1s1V5yVV+X
0Z8pGVCTyK7N0lKi8ya50+wl7pru/WY687iwZBhC44l28hWQPf9Wu9iXDgJ5dOsX
Qx/9kHnF6pHLU241LZd0UQSZmNnkbbfzXqKk+sqc1MehONqN9LhAwdaTkD0fuGuE
+bUGZ6v3Fys3CxMEZgOyEceKHtTdJ6hJJdo4qRQlO4Cg0GT0jTb34quEJ5ewgzwc
8TCHVqM7vH2nR+KjxsQpmc74TTIr4ysVMkfJhwI0qKy9njZLLBsxQzTxt654kQH8
EKG3qpIlNqYrKI4Aw2sG1dnMx9zyvqI3W1VgJ/IHjbvkBhpWVd9Gl3zYxB00I8DQ
Tu8so8JNPNC8rGzLQ9+xE7YOOpLJ14O4Bx1vSEngjUbp/XBTN3MkXN6tRmRCevzy
kL0UKuuccLI/VRKCKvXSYqqer2OWaCSXM0YlVro2ypHMCmzriQS3/LOFQtT6/i82
DbgY8dtIMulWMljWCGw8EAb1ql88cLDsvNIyXBHK9DkgkBUefDAPhF7K1IOat9j6
vMWp2idQQjDdnJx8wZAymTGbF3OGwaLbY8XX5Q+XSOx8Vh45PpEi7NDr+bygqJ8f
inNm/JyAQ4WsoQsoSDI+119mu+Hc5iHL4GA/gAuaJ8zTP9/Lt2FUBKmuDVSzQxd5
2ZmSGvw6NB8F2mj7BHb+Pb7SusGhjqNm5W/78NFbcJmNpr+zwOEJWkznJbJAL2yJ
vRDZmSx73/snPqpayXDt508zqlPVBg1Id6Ty40mDnvUtVp3l3uAeQGsYnkAq2TDC
nWaePDZtI8UYzSfRfzg5l8h/Jq829Ea6kFCfWmW5FHvRFIAwXE6hqtlgIVpRHCel
TwBUMC2WjXaUduICNFz0qVDtIcA3ir/v/V9L1qH3uwZxcGESDE2zOyd90jvV5Xx0
ZvrlMLBpqUDo2um3uqjuQ8zgNiB45mSolgXvvYo4nt9SG2F5pYs7DbpyVp7HtUdf
AYYU6b+n9Pxt4MUuyAcduXazYEwOts5uy0wGucboarhJq+pyGnUDSzzpjlsa+bne
u56lO6mrl8j/O/+dVZk1RrNc4a57AdkgXuNxjUUzZlQW25NiAOyLPAn1jxkSTQ3J
hdrrS5DrNaEcbAZwMaBRGRRPTTH+RlacWAsU8XXjTdLK5/u5pkV80AagXwN3WUk5
HGEVIBWb8vPKx7BTGBJcO6b2GLwJ7D4WrBXxbFOxduIHcwhKA19jY3Sz0iWVJBdD
Tmk5Pu8h9+OvvVlKKcgRq+UDlTGPcBPjmBqlxyhMBDOm4NQfaRvQ/LUo0QoqNISO
KB7ur+l/THqpu/d9uRdkiG4MdsaxPu/oaoCai1ZFbRtY/AufO5DeWk4MuEJXfRD6
7/ZFk1UjsrET1QwMRF3JhT3+7wAJcggESP2BFWkYUbNfUHzWkMjS21mzJlFBVe/f
v0WtXftP8Ah8rq/lxM/Fkr6NxWs2erQ7KgE3+Q3gHs0FI0PUvAGOHRXTkj4n4r4B
n5cnGxbU/BUaviG349WuhmpKm8ML2N+Z/cVHs3UQXoJ2Ufp3fBvbH4nCOcdX36H1
T4KvSWPV+XvXJZBD+CPp2KVC94gsNQA0I3v4G6m8Xx3HGJoqmssgo3i1xUt5k9G3
pFtozfnyoUWKBtPnsWptcu5lYvToSWG9D2tT62To6s/xKQYpqF2UTvMgy6UdrAHo
f/swGGFUGHroW4o/tTNtbc56NYH2qyaGXXNOwk1skTfNFGVfBLHo9U27iK9UtRx6
FI7yS+9QdEbeV5h2qMo8/y/3mRPiwhFw6jTrELUZ7JnPpd0EYD3DXazZ/FoWaI7v
nARg9SgEC9/GnWFm0vg3ep9vyCnMfpzL1dsy0CI/daqpikWVavIhB8KQwNyaKfNE
nUN54tkXzCwx+kAYJW+lVY/SjcPwOcCkGM0YCZoIJHdsWFZG9s+r7h08iHFixjJj
RlVlKGBhCW4+De1FyIAaBpYpX+9Th+vSHUDsnpXdukZcC8IyoTLhT0O1C5M7j7dq
zpt6K/Fg3Z+/bQZe+9nVk083TT/HA0b9eSOXZBZ7ydBIXgHnnCOubaZEk10KXYQk
TTGOT4QloZabQW8P9lzTEFsCWW65/+h8sv3y1smjhduo+aghkNft/h4zw7bAX/+G
UnKlLfT5zhf8gYvvtyiIOjCAkTM+dXMugGRr9jRquwgn9UqGN80Tr5KeyD3s2k2V
OIXd+lBSAedAliXEZqmSdUHBnlzkO3x0/d81zTFv4X/JGFJe+fmSu7dhJejEd4K5
5VzL83DGuJmerVL6wVg2gaOZqqjKQDRRqPldemXcw2KNjdMLdYTcbxjIqMiOj56g
WQ/uwrv7LqXV7uDCm4N0m5onKwQXFV6+mZhkCmQR+vPHk2O/Ik07bIERXVT89TeC
1BP9ZXdZ2qXbHUizC/LVBv59A0S5R3fP2qkJUhzSv3U8rjs0iPH40kOQRxhR55lS
2BGeSTi35S1lmEIX4TQwyRA9zIgikYmicOmMxpUCaC0OXHw8L7nyceuZzt6xyL9l
YGza8V/dwBcuWK1iIEQ6+6kYRByztRDiM1r0FxI9k1iysjM4Vq3TUK7n2ExZMBSM
TO6AYzCTabtw4yStwTYwFsMWFDmbpB8wofCYTom5MMT5aiGsAuf2/AII9w/GdHWi
/S+Yc9TcefS3deqkV0a3/V89F865wlVUgGVE99lwNLnl0Hjk1j/ixpusag+1EAzp
80+FG0jKMa6pyy4dRxrLWEoXkcoxLz7VMLL8Vec2iFSY48zsb5yFSjShSsi+xDjO
yIJo19GcPKkVWVP3fQiEnu+1LKGpE/XjfzY4FpPFO6wHID7BBzeD37le+vDKWk1X
LpyFehnBO2sUsb8SLp11jjVULfb1WTslZTfSQulszXXPV/RM5NGUOfIG4dHYQ4ks
ZKVCIlg2E0YZIL3GWALJ8SmVlYxw/ryyj2igDpIobTmWmuOMyETsHEPpyPLh8h1W
8s7Uxt3xsnt5m6ccOUCHDVjk3s8MKeuDSppDfs0zWZERd6ksbAjlgh+le647CFxk
b9w2B+vwHHCw6ukySocgotbvauuUU/WLTPHYtie9LyiRS10eWxHgoc9ehb5hYXtH
UEgaHvGv3s4uWD/59XlEtqpBmD1hjbfwNXKVyc2sNBZTkTzaPbRleg4syC+rK1Wp
dWcD9dcaGzdM3E9zTmD5hEm46pcM4KTU4muiPlWmcCYTdu0vRpWVd6VMeZ/bHf1g
3WhoyKpycnXdsVdYybTAxhn41yBKH+18uYPpnDT0JCvybMmPyX2/1cycOlLxx/MY
MkgLmhZDTjoL8R/nLhRaXyRNeWyoVvGo0f4xHhsLa6FKs5fsGjuW2BV/VvWVqKT8
hfLeWCTnPEzLm3TcCfA2M8bt2RW9QTUy7xHa6KT79U0qlnss2cbP3nAq7PeXwDga
cdCH6DsPAkUVzbjmUVEvzUWJeR5Hgsx5eXt3LY6/81ODliXjmycSrYnQKrrYMUCk
fHeLzOa6k3BlmfHzFijzKEheBf8hmskUcNzD8HtHaI0/UXfi0zHa6/fZM724ytZV
CJnJ/JhNhWc3pjgcLWCKN8bnP2EOhZSYejOc8EdkdKNxdqIfVpqlltaNZXcYEpsb
28WdmAn15Efpk1ToZMuo2tNEYaCkCVr9MzLRVz6M/tY7g8TCTgvKg4zC1Pr8DrHA
BIrMjcwJXS/uZDMm/6cDl45fGAbVJoznRQ2t9maPKehx+enxAsxdzg/U2rh5zC5G
AyVFBmK82GvoA5G/AOIV82a/6RPT2ipbuGWZtXOICE5goy9tbToT8Me6vIsdqcdz
T2VA6U8FUPEGbh/ou46+F/pgRtxhUBGD0oVuPBx4AnpScMScZxywIZT+CJdrvqBe
S6kRgw3EJSS3r4LNpYQxU+73Ddxs4LwfdrET7no9ZfrqCNc1OdgDXQQqIhjEJwXO
gnNOmBpqwoiwKoir5llz3WhlR3mB+dGxfHq+llRlbaoWC5s66kl52+wjzqsHo9yx
Ap3ja2ScAkgvXVHuesudZVYVQSwDK79w7GijvcnS2/LOl8+9/JB/1g+DQ1BxEBSB
/zeLiV1Dcp7kHPlCChIqYI78MeNCKtqdVF2xQNVVuKShjeqy5kySL6780Rzh99Aa
wU6fZxBcLPzIV3BBxej46dqMVJq736NCJ+S0fukPpEDFx9RLFV77T44pbAP/v4pE
oJGTqSDz0/flrWQaGnfFUTQo1+MgtlzZGLWFQt7Hb9t8CArlpjSwMpRdP9cUT2/u
WPDm9bbTUgso/g9KZPksGMM7uxl1dORkSjlmoDiE9WPpmn3BtoEoYKhm33KUVc+K
7k3PYGUIn0fFyF4uDYqiJ5ilsTslVEce2V0dG8TBFFEXMiINmA0wo69iTn+29wcN
`pragma protect end_protected
