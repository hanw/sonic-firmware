//                              -*- Mode: Verilog -*-
// Filename        : ast_monitor.sv
// Description     : AST monitor BFM code
// Author          : Han Wang
// Created On      : Wed Dec  7 10:13:36 2011
// Last Modified By: Han Wang
// Last Modified On: Wed Dec  7 10:13:36 2011
// Update Count    : 0
// Status          : Unknown, Use with caution!

module ast_monitor (/*AUTOARG*/ ) ;

   
   
endmodule // ast_monitor
